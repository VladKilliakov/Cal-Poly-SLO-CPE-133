`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ey4c1hSWFAc9TlRIPeZhYvsgM+KHspAXRgq+K4hohd7VE33CIDWoxnFS7PQIQEMwPkIpB8DuAujl
1muZ76ivmg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o7fas9htaCH9T4HZK69NxsUn3WiVnCd+rdI9/K1HcEIu5aJgOiaNVrtod5zEASSsZqWcILFcWzD6
Q1KbeR/smZdrsf6eWAhJPGQXp22BnBJZm6ZjKsERA+d55k5q3d0sXfntDtEU2DSo9aABzjUP0hml
UBXQTbGfhgDNar4MtH4=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TsUkDemS4KiOpFbeZOIlDP1mUsRTibCsco7q3Qwyst83/IQ7RDtOtowySsoZovC3nkhkf4PnX0+e
OPwHxr2ZGnqfxAC399x7USjTxU0Rf9QLaCredpadjZ5ZQ0Y9Vbd4HCruxx1PGIRxIs90bQrqgNaA
nUDuRMJoOpmjURFx+8U=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U+CsQMo65VtViMJoCx+2M1S9zH0yDaJhd+IdiISlvZpkaIv/QUmXuKMj5z4ZZ01IPEl4S8z6fGpU
SApnqAwPjC9pg8SUUFD3S/RQgJ2KDfP/G1EQzmxgEVjd6Yh4gs0iy8XfagFVIXPAfiXFTc94tQgp
QM5a0T/BTHFzGHT4HToQ+ROiJQREJFxtAC3FJYjLBF8F0DMJteveKi9HmeZbKsgRnuO7mRfJZiIN
shvfAJOa9LXV4Bz0JukzlYUC954RS4Hz64AKnVoh12JysVzDSMadwM2uCg5nTH+uBDb4OrukVcn4
1TlN/KInrqXV3i98VLx3/gOEmyNabA2qsPNlGQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Iku4d7TVaMR2gwLWQrFfKsFt+HQb8rRbd4/SZ5iNIqz92cSe3EQNd/7QsAOI5vuPmXx7TVbBHnxD
duV4ydry5rlbpSmDH7t80bEkUGvBpGlRQ9719CHvf/kfBLDkG786T7FyOXJmyVtWeiesViiObBBq
NU6c900t5gi4be4xYCZAYmX/hopxu1qFp0v2SkqOXLbQLMSJhR3UYMNuBYUCW5l7gEcPIGnxrLav
gdR+DpX35VrPWQe4l8ygETIcIxwYkOriXbwiu1wrBw09dAmqADfRzh9IptM7Fpvuf/sWKPq9hUB4
loPUN+1VTnxwPFBonTBI29Redyx3T3/QLmY+pQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mGVmJI+hgESYWxCBdO+QGXvKN8FJyfOII4LoQkjoPi5IbH38akbGTSbIZZuv9AfOQj7Z17t1Imws
PSUWg6HyJnWCX/lGvnU1zC2Qil2pzYGSEsOApmnC3q1U0O+/3gAO1orZUBE/L1kci5w+CheEcWgJ
0Tj8UqyGprBORI71NyFK4NfnBw8pKe0y0dN/hSJul9GRtNpUtoP+9ZgKcxzX288b0EhyFVdikDKA
Q1qv5xSo+4O1Rff2AZYwDvLnMxRQOa/QgcR3WEvrfn2zjDJdFLmpu5SqQb6vsKzNj9hgb94zjrfN
tWPUQOp6fxKZk3vt8EUhEtWivhx4z06A9WxHWA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432720)
`protect data_block
8z+VicQ2VsrqfpdBTqsGjSc7xOahzHK0GlCyv1Z3Tjs3fYH90wvzML/JcJCSamHZzTuUx+xMewYI
KY8wPXw/Y7dEe4UQQoKQ31zw+NE6+aE5tNnwnECp1zUpNeobvlITQyWNqvCcAJwJ2H/1rfeAI3RF
uDJftCt49OPewDCg7lwtE8+r1cFECFKY3thoaDRv5Wo4KXyQid3HVcUGrQ14BIkD7u4mesBzK7XM
R9RHwZroT89l1kg/B56NZ+a2pBvSlSaC8FiiuFoHMDvxr/BSDd3IAeFyetWJJJ9vpp2rXtfnPlLB
x1pRFnc8y1HnGDSYNKpjUBKK7khUz7T6iyPsw/mQl1Tk3FkSdZ0UD+v3cYdUSvkBUnTNad68Ty/O
La3pttWOns6BdqpIru06Zgu9XoHvvTqpe2KdUWXc1mJVLsIWsvP/LzDIy0Jsw8hG0wM4jYYVMt1j
6kLX7jwrKQvNAD4NYVJUGlTa1E8YDzGJ2Xm5tQMGuwfOPZquvQaPSeDEVX2bwhBRw6o1H1FOByKG
V04AsttEFu5h8TFwv0So2/d9bmpb2n2gjpOKa9OHrIKy8+HpljsFrdzXIdood2rOg0TMJE+y9eYt
1WzhcS40XfHELo822r8HC73LfMJBi/rLIvGEkYD7JXcI1Gz91e3h3dLLuT9CG+Cc6DiyHSLlsPG3
txbQy21TpopQ9uwG5tUjUnF0WOdsPvCXS5IrKjJB+8arIJFL69xYdFaeQk2fdy29S0/U9Ap3bKc7
CynN5szxQsK75Mh+8ABUqq0bhXSxW55w0sG/7N6ii8psAl4roSeZEhRya8xziX1YjwfPW31ctAmX
tZAdqq0Wf1fNDp65ApyVBKuiWGVNH7wUVHMr8trWVJVCsgk7XDNbfqczNmpsxQslWMvJ8Quu1CF+
iuLKfZatgxwcvuPu7zULJR/3RLGiiF2yEXcwLlEL821P0A4firGB6V1abZWmITxEXPs8PYuFWLHm
0/5wZOXzsdbSZ4EW1Lvff+4Lqy9h7Ntfwz/CpnJCmkeeU3qkDNEuxkJ0wOuh03216SV+nG1E8U/l
dIDILaFKV6PZdyXHsbklXp/2SXFu7KnMUTnQczuqRRRvDbnR34zBsrRr26ddtobcZVXYGMzixyeT
6nh0v5+b7e2qcUQSTPiIUaU7Phn2D7/YClJK1lfkQckbAE8LXWGNO+h1OKy6wjR4wGH6ykxiqEXP
mEYcV7wybyWzhwxAiljX6yC/G4hRpThgcOyNkobrlsvdkqPIhmgN3GxJV+fvlvcGlvW5PkGZ8H3V
RimpUeU2QtrwVyoH7QYunOZi3dsW0sJMEls2bteceemivqQmgNqw8XqNdaHPAQV4zgGrJ6mnILqk
qrAIKQI8iJJHWUKuSeIal+B/nIQyWSU92U0GrcVNsi5uvSm1mGoeyyz7DmSaOLyOBrrmf13IflQC
IdP+o5QOHSM5OlUFZPgfQRllTcCfWe6gt6zWhymaAXPLcTIOz/G5SWCCxJALIKwUYLUafQxQ+Hik
B0Wqzo+WJFcDdwdrXrzdSAM9agGe2FB1qrnKIXKG4w3Ecr045winuOL21sM6Ly3RKSIpZ2wEV8eq
wWXLOaVksg15LpV4GSgVDjg18258vaailUwj93XoveHxJV6tq2H9i3MNHcHRaBpw+NRSqthLzkvy
+ftT/T3Tnb1io7ItEr0egUJrQuo2Xd4JvEm0L7+ue5KTvYyZOBOYhN9Yoib/DlwrDihVF7yFWgKg
GPGlRaixiOHVoKHDftxOB90epVi6st2jjB38kYsNLvjRFqOi22NlDTrqv2qwOwNwC9ImgvMVl4HM
8sJWtiQNB17TD1RiTUhMSxdRCmNLV9MW+xzcVmHaP809S9PdWbJdTo/YtLc/xPe4jqI47pMaEZxo
D9R2tYHnWXfcqUOYtqWVtsO59l18ST+wby0Qqm5b1qeXhaumbRm7q++6Dp4gTKegUB2o8Xjm1vtM
kGuOWeHBfWp6GGElFYbELJkBHHPwXnVSAZu1ul9NNtp4Ccge89X32c54+z5nKpL2wbarWQihjM+U
tU4y1fsykrafYYeEkAQUcb8XQFinYL6xcAJLyfop7LF0dYVZ8U9Qt41a+dfhSBxaJVWd5Fu7shqs
NNtO9JWdtMyq1EyfOjAXos2p0jMhXsfC+dU2aqhO84YihAus6XPE76b2kbQd0f8jr2YjzJpVdVAJ
70c4Zc0ib8e0iMpYQGTjs/xnHlt1NMvQT+XsBjATufX9ZPyIsJFjCFRuREKNAQKs1sSQyCr1S6qh
sMZBmIKHysBkvxkHrN6MJ4uplvsMzKLwJyb98jE7+X41CmYmQPmJnEDA6isA/ReG+YidsCiK7OLM
zrbaWf1BBnhzeUZ4eVOf7GcisB/6EMkgpeQIm9I8UNT8KhBpoGuSk8ifYS/5I/V0+gZax1IVxAZP
KSOGatnVSlfSM5BC7TfYR+cyNOEwNqbSZ8VLlDi0yZrSilFmj0M3Cxf+OhJmFkDi0Orywgoor+iK
LqM9C1PPTkl/4EbtKfDqg7CpwbCN/X9f7n5VPjRBEEJ3uCOgfGBT8j1hdmXuujMWvtBSXTDsm8dL
k3nPNq06AFbR18F/5TO/wZJt+BKw0b2+66UOTR4+eYBu0YbpBQQ2CZgevkUGUDmPnVxP0zTRC4Cr
FIan9VWm4LJ3gwpGdbKbOrhAyJRhmMG2OQdtat0qgaSGcCdaKVFfiU1Ik/bXZrCDzHTBeqPQgr1v
UBxb/whRp08Fjw3c7wEwwpuN9Y7NjxI8HmMOr4I+DPmyyVMLMACSm/dD2l675+AVwqhw1RLvDdR0
EsGwzwAM66HRWWdAgEZ8cq7ubmzHXJ19glGCqTWZnRKiqzUqU1vT1XkxVF1rWlCE578iEmeGhYGs
+CCE9SxjpU9dwZwS69aTDI/SRRZGDR46CGdqkxa76Syx3QMv62qtC8a4pPJtc1lk93aVkMOiV4UB
mkRTsoAHA1DV2gIPrJhHdylwj/v+CqN7zWXAmlgVIgz8LEnooQyGTfsmLTB/F1Wu1ipFp6zvJCJj
t4Mj6Ft3qujW9putQwVI+sSxVfp+16M3CANwbYExCtu/54A0gh+rdXbE0ssq8jwg3u5dduplOHIL
YN6AbYqVHTqwmTd+vRVVADc1ADKleRQ0QMDlTPXbknBC7Ym8321IJg3y2jpXRiInk0zARdWuiVHA
iogvjAqgxaw2vxPBvsFZc/8HYtGhzYdht8TJRDyOilNaXQxqCU3mIKsH+RxIXUAioYtMO4PTsD76
gyZE74ow+mabJ6x33kjWziDotQHHsLxoHa0+w5rdUccRyH75KRyrL8zRsEQZ7sr6FQP3SAk+uv8t
GB99Sz8OY1f1R8bSLqmrTB7JrYbl0EYj5aLOGeZD8wW3AEYzn31JG45ksJ3CoB/7HZYtz+kpJcyi
byg51RwTVWvzzb9+czLQwo6oCw2gc5vcmNScPqimYRBOyVPkYhBzCdhrrC0qKDdfYkw9oXOt5mKR
2iaNMZ29yKvL3Vm7UUjWkqR9q7BvEz1d3uLqOQ6XaKmjUnzKQJe9ST+4DGYTgLgkNjwg2+eqQVnL
2Yh6JM11rX0KRuBtmkOrTWPJ5HfnsgQGIABCi2oqjmfV2xvLF3WKyi0wuChSHW1N6cA3qWPKXE40
pUL4s2sl1s5m1tPml582YrXjHzKEA1V0dWPxgA76wC/VvqT/FhdcY5Sa62Dz4piIs911xEB0NA0B
onXEJJyvuOsT+i1b9ciatRex2XkRyxrsU722CIFxIrBW5tfppuvfM3X0PrBxu3JBYQki2AqGyfOU
EMcqUefW12NAOm3bYfvgd9L2BzGES1G6BP8+TYDeIbNaVucpp1cWkT2JBizTCyr+Q2X7tPiCUN9p
McMBxfVnnbQAavEuoXnhTF/akTStcezo8cOIQM+ChVIAZdY9jGQEoouzG8ThCVxhnQr5JEJmhew8
exH+YRRH4zCWQb4VDD8GCKe3kMVvdVKIG8jwZAViJglc4Hfo8lgT6QRP3zI9KVm3DEsF5cIme0lU
LKc1Mp7H6vhW30rZ+fWCpYXAecg8c94HdIX14hhuvdB9KvxsxytiFF23+5XL8NdQ1R4dDzPFCiVB
pkbhlIqpbvXJJ4+RLodolitoaWH7FWO0PM2xRprbRKk+zAM2lXWxHMhhXGEJlA9SfcJpkz1fB5g+
i98rGAhet+Iqa5f1UxaqVW0dCuVkKfJL5vHAj0ZU+lcAy7q86j9lDnwQJTjtJ0SqgpkwMPHvFgp3
GRGGUcigI8P5F79VPfQcNjkLQr6D4ZyMINLEslYW5lLbIaQOoX9VziaLehdUtZIXXTSqE/bFCckU
fncSaVSTQskhoNSukH5OG3oSv7218idPXRHofj8vBjawDowp1Lzb4hrO7YtY+UbbgU9DUH5feGCS
s4Z6aD1Ij9BrtNYS6f78Y3EhOeVMq4cFtU7/rDIaZ+LEVYDjWNVjACAjExSRiiPQtHFVZwK9wy9W
+6X0s5ZU6pReuivbcEjobTyQ9GTm3+tZBRF1nl+ZDlkrR4Dh8c3Q2j3SLY6Xov1aqU2oK1NwcPHj
pobaMFxiITtYJz86nAumUaUbUe9r2WawXAXre+mxtJPJ/SWE3V5Ooyi7HEUJBHb6B+Ml14tLOXHL
jnphpOgIvqth7Zg3o095T7VzeZwWFJMvnBqtxJd8ktCdk+/LYz99QBCylHOy+iOD2ylKMAcxmBhi
rIdwlMV9j/RGMxlCMCSmLCrKOjfNVWM2Tmx6PC0GeXQjzUlMjiOc3rQ27cBOOZmWcb44iZ/t4L8s
F9Pp32Dh9F/LUjRMnNx+SPHrX2YtQ17nkqaL3lAkoCf2fI+mjMswNzmPRrm2Dyb7cM7s1OUpphBi
jx8SLU+vvQYLo5CtlDhQpdIW9ShScdbHqhX2/di9dH9TV/ZDSiBkLX58Fx7+ISJ4492SISuNb3S5
nCBHWwz/NJdopJc1TQzmWWUUE+BhFwqNL9EXuKsnhQnulMHi0ehJvtwxWozmRoKbX8I5RbHFyYIk
SRmGytzhpkEu5V1JVXWmrBhAmNFArEg8qvajRRJzZz916l2uXiepnKVGJ1stcZWYG6tt960s0mS2
HdUS3ESJkO04jBk/Cdj1utnOOsQQoG6cfzB/VpE9hBOtJ2PDCFu8Fzzp2DQfeuuStGsoQsa+N8HJ
ZjQGKJRtLb+3ScAEaZjOmASWy9teyQ+YvDu5JnBbVmE+jj/wahDQYP/S2UahhnyM2JekNdPimrl6
lC0zcQ8GYGkXzzZolG/pYxUHRSuWUfBe5j1/iG26kLxX5uXwUneUXs4bbVcgCm5z7eGJFVMe6aG1
Rzt2kjs4DJs/qPzmLJYzbh6SV1E35I5+4yBDHGQZgxgou/STCqffsgq0vG9gs8aRL3ky5Momkskk
2Fg4lp7blP4ejFUpYh2OyrCGmQxH8xFvJxs/MjSO2cIYvDhKbyzSIdPJli2/ptPl9p1E2v49bBRi
GA7x+XS1w0v5Ku65A7aL4ZmOc3A9hNlmqNnuLSyUtX1EqPM6/2M1QDDakIdayuQRCInyv2jbjDM3
7JO8vy6PNw//ITaqdSbJiYhTXC7LN1qVrXHdr6hlVloFE5CSPAI8gezVhnJSzd4UwoEWTPoms5OE
Zb9B1jnl4qB2IdRrTCkG6EKg5ex2w83n1IUIt1L3hQLmeJyvdENQPaz6pGAnXklwb5uFvrJWY935
W0T0SPvvZgS8eBnP3B4mByQkzH9VXOiOIlMwYuWxZLkWssYYzpBCwrpCrS02Ngg9ORfUfwtcGZnt
nfsml9og179Ft7YCr77ouLN4NVdlzRyTs76OY/2F5g3SSVB0OFP/jBJ3jtTpVLMpZ5ssCxtqjeNc
PLgG1mPqtZSAqeWlifjg9+kKIH4Pm6ZBj3uBBiopiwGI1NNZnLCgDHwn0JSgxytYkJ75GP60ToHR
zOzbgZx0N8v8cNS7RnRGdQUDt007dHhg0628uhcvn0sr8mNiBIgXkK/cbCN7JISNvjzzl5+6cPH9
EAOqyVHlO8Tn3UCU7zAfgLSzH/yDLgzYiaZ2nbriNqwJ9xbtM1B+e0ySW/jTo9ETZaqub2Env6ET
msuzNj3VpYDcfIOdgKzCve93/ejVy1se4fKRlROGESintnXbXjRNfN9vNm+8q517DhRdSOt+UMjA
3gc1IrQPBwxMngeXkJKKMRqVo2u5nXBq242y9E4fUzg9p9CXSKypn6jc3PS5LSIClPak9ZjkhSK2
gCeRCAT9TuOdGaa5waP2sRBg6g7iiyqKD8WLtoipakIHjPko7Ha8DAAtJaBmECPOJWNtZ7NZqFJ8
taTafWwcHfi0KFNGo6tGL63KyxoR/k1EZPrvjKGZSNJJExP3YH2YU6RPRc+lZOp/1NwdTC1brD88
u4jtkYywuoDpE/XCNQhLZLW3i1ipxinDmFeIZQhalEsgx58HnzwbuL6vFPOAirbel+6xRnR33F4T
2yKspuf4tj5xdRKOW4YMXvHR4HB2W7OFdjvMiy0lv8z5/4aBOmuY0BrMgTYBS2690mrfdVURA9C4
eDIOqQbEMzMr+GgJvZuM367Jj1pi7OzF5ExcTUXr6oVJ/ANqVEVTIri5VOhSUnNQ72DsXYXRtOiM
uBmEAhVMInZcNE5Rnwhb23YAUYIZPN9rcQpKMcyRMF3YUDKbakqr8QVj6VL8y4LPJCyz3lo2XRMd
ZoDJuMa+EJ751BiPjSmnRRcZCmzRLM72C+KwMawvBzx3hf525v4Cnw2ZZpedmGDDXJgFNWzfjMem
09n8QpdB9AcpBXfGOoc9CKdWnOOoQQ2LdCYqDBwaUe7DuGbskG6NNh6M4UJyfNEsGv+otu5x0FgB
mwMHOf651Y7QtjRR1cRFaRLTxH7Iz/g4CMS3/l/hULkefQNmWjslC/GVX8W4q1R9e3sR3dUXlfF6
XiyOf7xnszSL8Fh3jz6u/DXeKetvpI29tUVJOy/YknwKKfa23v5i4GfSguE+u/1l9fWLlzkkbBRN
Ej1Iar2BywXaz+FWrt8NRCPhnAsSXIWSADCWbpHvE8l5fGgFLWD0EI2rUuNHXrvXyHFWHdSFY6X/
Y2cTkX2nzEFrK9QEktU68SIza1fePUVTUUXe1cSB2rilQRV1pTUbr/pvqDen4cGTUMEaD1KuDUWG
ZRqxdtbC1c7C50XNcZq1K+CkQQDyq7/y5k7NtWtGpWa4ECum9DmAHjW6JTw8BjF6TDMpCUBYvBwK
KRdwCJA6Js/5v8oJXeGgqBog+QmkGkTrs9z9YjbkV4opGrdYUurkgB7OPgmy64OmR6U1yV2wnsVL
/75D4BZRZJYFBLKhgrQtm2VQMq1HkLi1K+ltjIOUpMP15ot2m73zbWwNRkvAEcNhSyu90MEyrvIl
2eMQnOPMI+psc6pmO6PPNQHCXGmV8fdmz8d1f71gaLCbL9WPSzkU+1H2ApVLLLevbII/P1lSBjQ/
BaaTczJ9b6y3t5qaCJ1k/dNWYu4iGzRSj4NKcojvxlg2uYD6BzyxRAtsULaLyu98CnLGbgq6kFoM
s/voonuITrCbpJGjh/E6hpS949LI+moc/DE4YtuepVcHxoHyOc1cdXyv7QQLGFn6SU9uchUFoXzf
enmwDc+Gcs+c3irwrbWsnVcUYcs7pUQpeQxlQd05LWAg7b95QCYK/6mgfn3YLDbPRhOkPA9f3SCp
FWMBM5rqZm/IOZcRGzNwMjyELwQVmw4P2Gp74AULGs/V6M5L6IOwOeUe+qiVQeTYvCh95N9B173o
lkuge/YtRjxYAlArPVd5TAsetrbbDh9mq8HJ0/ebENjwui9VPxEBlYKP9FkPHo3ZC75pmCVTuDnG
E7qfvexSOttPQfmOZqvvCpsrtBdSaFq3ZoG0YzG+kYlTyWkghBLKJ/Jcm2o6OV6tYya/uHLWSOmo
HJoYxEZtTaFYCln3EE4QzDGOriG6BpOl0iqaP1h8WZ2obM0IPxfVy/G8lgWPSKaTv66pZpD7TMPM
hWDhcWeQF2/5uUFLsrZvVjqOSAjYTStEVhOwE5yeL8n2CBo4vkDaE5Pixdn6ooNEZeShYV1nXlbX
1vznM+QWD+khBCpbiRWVZ2JsATyt0DLV9zepsIfxd2lqSBonaX4GfefRYSj+3HchOtj0hrkHBUyD
ux0EhpoAD+qE2sZKccDA9EZOPsTN5K1ETLUOX60Weitjiojj0LZQURGx37DboFsf8AbSBXG7GSQx
rR+dNIe0k7s4k9p0msWN17V06Ghr3EZ4cmhNpczVMaBOXKBQI0uHxzJPkXEjL1UISLTLYnE+Rwu+
IHWB5Qf1xnMZsluTaYu5X0AlJC2MBh1Z18fbpbAWLPfx0JPqMcCi8hlHXQOPh4/Q8eKhvUuHIXmm
WrHErsq4OwyUNdi6BAuYbfxYVWt+0wbAcAlTjbbLkvdT/BgEj4kfzJI75nL/uiy9c67ign3xXDIX
haykuaIYsCQvLZpzNlyHBWfPVuXPstGvvH9/Y/e4ep1/6W5TZuF/LAyc2aZStbsWFnbeXw5Q3gFj
zC65xUcvxRVrmGY8m2aBk9Sb/dAS3hn1Maqgljzw0D1N7+kBCZevSxjnWjFBoxTRFfSZbZNFm6DL
wccxVQ5vPw/AEgBLHPzEKtysYo6PVT3BSPdgwAR8Rv4zlJp7sdRR420oS8SNKtnKs0wiOCYEP2Qv
I7h5aldN7bmX1J1BouwJbsbLBng7FFIutVYbQO+ErFPgJR7j0ECIvLnGL1DlKQHRvUkpnZSwhO37
tSj9HK+QCZ4O9AfpBVuGyim7XFDIW/nVXSaiLcV3KpEehhbHZcc0HESq3b5wPdwPQ1OogQPrVxwh
7ne13VCgncfsd1Ax6iDlAcubN/UEjK6DHlPdwjigqqPIAJ32mFFCbUWZVzj4LjHnT7BuT0/hJ/Wr
LY6F2fUcpXlPt7oaESAG1Y/+3Igdkkc97qLykzuLCz7sYl5mGZ5a5kqhlYi/lp2stpB15H35iCQM
kgCINf9q8LfuWRMJjDLsXdtWDi6yO/OAruVC3cTKOZpTPnmwPtGZSa1b1iet+Xsd70GJJlnj8W+v
8xt1RZ5vvMMczDAcCs+oaEmSvQ0/FbH4hcpBAm6SA43JWCeJqc/KQrgSRJ8xJPX6hzI4648e2FZb
5fO0oaxd/RrTwNgdYyZwc9K4vLln9M1sMHt/NOj8TwiXkHIHzgrvKHA0Bkh1GBsoTVAyng3SQ1e0
AbDZG5SSoQhEnLruPQPdX2WAtUzzbcM3HkJvk1WB92tSr4v4E8Gz+MJBHbph8VACVHnsCNPSsIZf
Ufo9iKAskf6TIWsPcy9SrWVeXqfDX4P71Dz8V5x6HKJOIbM2Xz0PluwPEncL0eQiuxTKZi8vmk6k
MRNb+f9AwpBF2+4/RKYZ3iaAWKyrmPHIwQ/hE9K+WG/HtAtwzH7nqnd0qbE5FYZEq1WKxCddsURW
RrR1r01Do7pOwIs7sc/9ekZ2X1O9mTaAn4r1jhY4gSsdVUkEFFbVfyyPYh65BOJZp1x9gOXgalSD
rSL2Np9cHFC9luzUx9uzCAaRXO716edyUYV+nOSGhQg8ljGtFDC8AAGt8FXDkZXIsa79+O7tPJeb
FRIKiy/KTietcMcUaRAm69FKhykEyry5zRx0elO+B4YxqAQtmm56OuzuZwHEMom06vZuisBA39Sk
PEOdiwtNIDLal0s+8Cl6TT8WM8axoKj8snvYcdGZ0kZfR9HSifLZCrhO0pMn90BLtxsgSS+yoapU
5TZXRbmaXLoWmnyHGW4O68ldA2srr2EhwiyIOohu4j/RKNYT+9KGJvSE1BmKiwkrWkWEKFVS6xAC
KlfVDe+1hMUtQbZKRgl+YLb0lPFHo/iCHrn6GPm3venRrAeIdxvsvpfQMy6VMAkQ4ZyS+rxfN38n
PNf7U0ngII74RimRW+kzCvon4Qbr4XNGqV9p90FSklMFb1f/8wS+ta9UFYLrIiniqCxWIf5fZm/a
lZxCc76RN2XG6+csltZitNI/WKAZscDLIyb617QCt/h7oMVPEnhR1Ushw03XM9gx3EQ4nzcZXYCd
XJgdOj46JqkqO5cN1sJUscTIIQ33f9UkD5jV8VoBacNHHXRI81uqpC8voDzcBy1llvQJg77Er3aB
3HwQhXtWJhya+0W7gXP9VUtr1+y7zJ/uuQVdQgTX73Djdv7ng6rVhI2BPN9At90cFeyOkVMXlkTF
hZ6O/ad8+SE0UJWkXP2/vOLLNZWcZ9ABg3E3QaVGHHM6wV1c7kWqQBsmQ56hFY8AnsKp/haO/2Ib
0jisSumwc4LIRQlpBvGmBYsffQkeuTJpePvggdw/hkpwSiXCgwV/9bqW9ryAa5hhKvof8CgrSn7g
3soX/w6r6gsBHhGJJcrB0Uoa1aOhZe4G5y8tX4wOd7AM9RzTbe1JDTgE6FJqTQ8JQ8F8cfC1lNyZ
wyqJiFcCZBwCvXTQiH7aQJSOcsIO5lP+zjIAEn5T/oaFUsApSlyI41ud7CQgaOGDAHZXRgkD43vM
oyKpXmUiNl9OIIR6Di/I87gLmSeg9O56gvI/dWk4Crsz6KfXqcGZmhMbMrwehUh5fLys5aVBfHqe
Ri71aVRRxsxAeGPPgKXHyP5Vxgl8tZ3h13vcqn34oAXhXrvqYZCfjzXvnxO0C7v80gtVt8Zw5wVF
8RGQVo4bg7JQHZ3jgQKOrTWj88Wu9Cz0X0BHT7hxwJOEfpZ4tyN6Nr4+scVxJQia0ekuE42LFRvl
4uc6w+bIml8grbj/PJ/ReyVaXQRwRp6BuDXP3TcijPhtQ+Esw/1W6DDnVSIHUrwPuxAitsS7rgQG
bOL6tNhLfk4UX3MZgBje1h0PNVNMfXf0rRveK9anZjSuTTX3nvf6GsDtV4PPPyI5/HKysBZMZLJg
fuUYFKTmz4VlPK4S/n9c3uOTYqraI51wffng13PqwVcpNAXqIY23e6WhJLBI1l3kbrgJJqYULypI
yrey+LY1sc2FyW73hW+KNY1IWQUD82YPwg6QfReLA8jfMkD7Lc0zv2JcYWv7qe7lpKR1xmP0jdhS
8eOHrIawaTLqImR4GzNFsUWOFaeV5lw2b+nsolquSDYPX+q2AIkBm9wI/JY+lATzO0RkuXU/aehq
zbkxO54LfwS4WB36SD4iw1Zd+KIIkWszLWWO9x8joulTSkaaj0V2oP43PyGsPAp1+N7DLgI9/0BY
xckkEC1GYhTHbTdZha9g5jNUKFq+F989/wGcB2WW5rxD+y3vVMWjjX/b5AHTb+JvZ0J86lGayvX0
uGllejGLe+GycWuLCwytrrFQ824H1ilSiVYt8PbMOb3YPt37C+b4uhq7KtuHyqhZJHjsQQNeUw7n
H34hrcsxRWAizvZQrsJH1wJHE4Y1LGKre9kVi3ogdfjVOz6AQSpAU1G97b+c5LZV5lzGZo+Zk37q
ABDn/03+W7P2WD8PY9p4s09aZAQInS7mTya+DchHvavDvJG6Xks+WU6V/b2fm9L+7gTahp6OaeFj
h+8PHhuSIcG+/a8SAVId/05SBgyfwxU1sjIixxEO0FH5Dp5tnp8mChHf17Z645KqkOGXy0cQwL07
C9Wet/5GlyVJU+c2X0Kl+8iTdzabRb5TjVRbWLAEpWlTEYH2l5yxcYvXHCqnDWooO7UVEIvySodl
UYHkssEOwbNVkQyd/uwempsMIH/Utu3pBNl2ZQHroGL5TAVnAzD0W4p0qWKfnu8GFwb1/yVyJvIv
w+TEvCOpshiaTlo+erlRElWPM3HcRA7IwAX4m42llOadJ6DQCVJweucttgLFjP3w3BMloT1uEd9p
Gbq25nXamLdCPaMOk9F03O8/OfWYZtoSyHQphV6OXpQPH7eo43asSfsK6r93azo8G2wa6+PupLxa
GhCGbKte33qr4E05qyfW+Xn+ro5u5bHzQBFTYnXDVGL1x6eKWOffVSIjpAlER8syNm025aZB438Z
ykTIWnd4JbaDKRLplpM+nvZ3tiRlonHqpg7yW44tpD+qqRLCNp5XUHzJsfcXSqbA3DuIcPHYddC4
E5kdSUrlCtzz8F+AHbggX1AUBriJEpt9RvKZ7HAolku6sX17NOXQ+gso1iUDM5cTgWywlgmJdRk4
HOCSeHzzQ4jGymlUeOzMFym5WTbMm54E89k+p9q9YI1EP327c8oE6TGeVjhm/l3a4rPh4ItMeCvc
8o/RbZ7KlyH6wdV0KuE1+nApEc4EnpBYaJDOW69vu92oqsvRLkqRgR5ffBd8iio7s99eAYB0wX8h
wyk7nVslE2pAKRyZ3gfFrTcXET3DDs4tCdgEs/EAv7whpkJZYyn24/Tu4q6Y26YBVQmENBu7w85s
q1JXKaWzfUYoFa0814NV0sHJjyhuvRscl6pUza1qkRnEwoCynadCO/XVt+uJAclO2beqqHkOd+ce
ORoUBMsTmO+eDcCJjZ2GCvebmIqtMyKJ8vXbFIV4kHqVSTY56PhWNJL8FrO3RLsdV1+wlhfaNOxx
DxLUIANGiCy5aq7mYxcKu/+ipM/72MnNHzh/lSeDe6Kwx4NuslzAKpzX7lGHOjtH9OZrBoL/7JhD
MJjqKTnvIFDfUKtypu38YzlbxdKDj5M+OLuZ6AFR3aYJPXKIsU7Ju3HlzDg1xI1B1gR9ITjWFu0f
pBdiBZ2qGwoBji95xiuPGqQSZml9oPjTOXF1Z7nZPsicrfLbNIuWQV1WJpxKPALGJayulBWo9KgE
EISIZGUhCn3cIUbdKqqOlfx9zHfOkbBH6YhNH8ash9gSzFyy43Fl+Pew2a1js2iUSPuG2eQtYiW4
HDRAA8y7cIKWIEYsXSZuN0HqTR10VV5Sp1K6TOfgE/4Q1DzWjgFIzXYqTBpla2PJBKLzIoCJbggJ
0nsc1mdDzZ2ZETCeQl0Tz4ecRfwqlUu789VQ1QnETKlawTZMkmqBGiBjXlfmneMudcTWQt/xvvoo
Q9B/g34/zCva8KKPAGEpyynZGUwyISEm2BecJM6KuDIlZhDT7n5Gdz8cIapDZibfXDIhST+qJAim
thrOYvexe/OiliRw/yn6UzkEESIek0Ld4Hbx9Bt01mrT+zPL74U2laMpd9X+p+I/bXA9YLh8Iuk1
eDQQV9J1zMEyUXz0FUrSGzoaVS77ySd6A1uXuYjC1iGiX8ZnZVVYLtEDgcS/e1GFhb+6D4OlYLDt
kbaeBWYeKxl/EpwU7nGKQxuqbuj7q/RUuXTHN3PcG+ODor+o51gozH1bkzWWFw6ovhERJP+IHWLt
/Q7JIWfGOnyCm6tUsDr7Zle/QebLjRYAygl5+Hwt9cIe/Xr27XcXM/ybE99073sL6qlCYP+ZB2zT
DfJXpwgHfaX3VVzh118tQGkdhghkisEmxXvSgXDJm1+1S66Wzj8sQJYeT7Y+1Qd+fYKqUirxFCvV
E0Ty99YdubS7EDkhEy/EuhyPdL9eubedQdAUI0YoBshEU5pa6CobTa5/5r3RPGdwlZNlEZcrkNCA
WlzLaGhl/YPUsn5gIwp53sicuAvjIb+TXbcTez4DJ1ebEnzd5UQTd9ObDJdw+Vj5+SZoCnS1OsJv
fSepX8w3N3s2d2kvGj37PcTSea90vam5LhFahlcNfMvnGM/8PRbtNQmkYgP6kuGl25slIho0ZwpM
wZpsovFHB0DZzuAKMSv/atgSnY14iY9QDQ8yUXSmH6iJ3uTQYSVum4h889KS/8kQVnTFPPJdCqsX
YJDFAmcUm1ZNz4j4ISAARfF24r9+A4RCVilkBs8p32kO2or+DuSNnnji8fGuCEynH+bqBX/PrE/P
K4H8Jr/LXiONOjEZVAEc6eP/e3rNXrpsSL/L475XgEKqwvVgWRRF14vkmSx6250YkoJx/XytUYv/
zvjN9CJKstq+KCzERSo2vzFb7IZ+hnTvsta5pvtN9zQ84t9xtnS0FLYmhCe5m8b9K/CO0FJ1mD57
cWehPv6vdzjFsKLohi/tHvOYteYBgqE9uoIEoyPTP/KYpBIhVi9qH3XPFDh4xLR2hRhR/1YcGzod
hsy1lyqrF/HkqZxybDTqDviij4HV1rZn7NXQ1f2WtZfMpGu6Z3HiZexaKem6SSODms/WGbCpWREJ
lEmc6OrYnnVvG+JEFG2+Aa2Z5GuX9TPniHqACyXAjon54Vx/yb1xzVZ6HXHX6lTHWmNf8Qa6X/86
kp99ZUjL/esaMQJ6d85LkwMH4PVoRhS4/9JZ5pu1rD3LAsFbvkgdaPNF+UENjVuRNhl/dO4GU5Kd
MO60gRYEZ1QFaMWhlez91nK3rz/bfpDboS6XiK5hsHXd5oq17yIh086S9UEjKn5IJi2NeTumOPMG
dK0J5eIADyT0rbOmGYUqZ4OzqodbWat+hsNn+Ef55IEkSfJPTLrc4f2dQj8fnVjsgafUCgt9dQ7Z
qFzioRvWvhfDNBiCvfS1jjtzYBMG4CESvJcclldZyQ9jeV85zYc+SQL7nhNa0kU73mELP9FKJ+Vs
F8SLTzUxsEepm31ViP6WmyJh2Z3zNyy6miWpe6iN05a7Uf5Y5RW+QbwRjJjFjNy/0KSDRJZ8K+6P
uCsQ9d9HuQSyYimkq7aNhRM9uypmWsKnXESm2xapraBnttXilrElIYs+Ckply4w6xoOW65zyeriM
XYT3DRbg9pXEHCs/AZJW1ekvUbHfl3ke6TpuX6a3GR2vSeoNDsFSYt9aaSuAp4BlMLcLqR/kEK9K
+sg86zOAsVmwUM1dhMhnd7Zvd6+KGFBOYZLr0jAxP3BLaX7EGX0w5fVIDAmLjN/vU2d51NG+i3xu
HKYTBqWlSdutaM0aT9Tjf1bysaVY94ZdA0CAnxPYlPDREUrHGoEBDEv5IWwv6FTIm71atwz6IF5L
B3uLso1YRbq9yRM/Vg3rCmmB/QwLkWMNCUCDE0bHkKr6KhsbBbQfq0o7vkX3hl3B5feuPDeG20Iq
kretIJLLdUgtCEWT998zPKve8441TwFjWohqs4cZfeHjUcjb/bUvqkwCRWXSBGqmMln4f8NzFLAg
QXm8gGxWP7zcGO1PSM4YpVEehtNDfVnFfTgXa1zvVekd6kM0kuPS6KJzsSHG3SPF0bHnEXo+tQol
22RcSPGyG0mrOkQxnH/rEjuOhCfJXsICJppFkmjDmiU96rJ9Mx7DluMhjOCKMCFV2JHYGLU4VaNJ
eWT6TP3ndK/G1lqk7ZnBrqR5R5fpCT9PsD7EQH71wmHHjhSpPHrpleBFeMcrVRQcbKQZrrjhFHY9
JQ52EWcszZ60y6ULQ43e+x1yHX7+rjOgxyn46E285f+FvicpMABl8M26kjvXwj1FthK3fImenYIK
ViFc8RBzwpuf6pfv59DkzBVb0VA9FU2RKWQyzb2RI5igkvejIE21Bjsqc/Y+QB4LcBH/vmL8wIKJ
w67q6u47D/5eouhgX21131xJT6HpSkTa8J7GezyF3yBf3ooiAtw+jsSljsUgFsutDafnjQrNKRxG
Izryin8b4/JyEVdW1XV/kkrfpSPHE1HLlVUoreCAFTuXJpl+dukRPTuXM2ITgX7rNRDX9JYuKeTX
9k5QpTahdh33ejepJD6nFH12CVZ9Lpk+t476nT0oi9iHnlINNn3RS8re/bkOAz60PZR7JlgyH0S7
cEFYKz0+TMWP6hHlbFvCDDtsiTxYjRabkn/NkUeVLjjw1c5k/2dQXiVhlPtHiiTUR09dSvvKxgEb
VffG2k4bYOlIxvlfhSRJ0wfZ9NlR0kHYZAM+hQn1MriKjxb1vAIKTixEOEXDieC93JH8oOHBS2Ro
QdxWXV7HA6FTdJobP5Ij7eL2YmJELj39MLb47VD7t8tW8h6btfeGdMkyht+VlIflx2ZmKojVUrkn
nEsAWluvPmGH8llA3CkZwUJmb87HXRyT8KMZRyiBNi/6Gn5eER/1J3QkbBZudL4s7wKqfH5AJG1c
1gIYucDH/UJarNxlwwUN88/+CSHDQkdjBPzl8cPWGkPuv+Z02kV6HF3YtSbByyrpGjeGdc9V5IOK
VxezjFZUCv+VscSxqRvYh03hUTnllZ8W5vO9VelpPuMiR4FXz44lcJIpiCju33+ZiVdtSadyyFoE
BEvbs4FJdhICTksDuD+j6wVep8W9ZHU/zt9TVwjBawAwg4l1iLRXcqZERmgyD+63V+JNgSQ4DRwX
mV4B0CZ5laPPzc/lXlYlGdY10wVek5C0kpIL9l+dXbDf1OrZ+c/rriDgc6NrF6tvASXbOqxdi3/H
vrsuNPcc6i1tG5zDnPFIY31bvBgncnhzR7qHmr/I34hf11TPUQ/LHdYStKvm+RfKoxrbvAN5A/zS
s01lTVRI7pWXUZ5CMDEiO8nZ1LlBgzuy12ifWBMSGGy22pbkanjjC3ARH86jIHrqsr7Pn56994a1
Q9TnFurXtjrTcpL4zt1Hs2cpKhVS51JK6RJPaUkjh5jFT/sLdHVf6wmudsHcLnmlUS5ITT0HrHTY
tyGJ2N/tBekLrSFdyv+QtmM5f8RhczGByDI9D9NtUKVGxW1rvUs5FSUEpIVxQynbICJyHBe4+DF9
HCuJswcmRyI7L+7JaAiLnlMqDpiplQUFP8SEvZyb94V6tEHAF+JR7dw+e6Daf7i4d14gqi5sN7dv
HLb2+OBBTNuyjRvrtHUGvpGs1vELUEpN51WQKfwPGwBT1bE+rhFGlNP90TYcfrbYE8LY3s2VBUfU
kddDu8T/pnEii9UWMk32LvqqJyiZXqbFEQDLsAY3NgmiZhzq6Rief7syDpr9/GjdZJyE4uJqa7sb
HrO8c2ANPtuiQZuD+LRWZoSJed0E6WlUUPZD5VS1CURxWQ9mk+0B0hasiP/iEzi3TAb++bahrPGh
WhoiYIwuu+9kSFu0sCM/eVbEQc+pa7mG3MdK9VKK8jeY/0iUGFJjoci4i7UVXgiQQ195YTj+EFlJ
Hn3QlksrGNS4bZFYSMEjd/jR1JKrckW++C2gwBBnixQRW96tpFCtHp36rxOW5pGl2P3St8KItKgp
652bDYA0Bz+DMy0htCllQTf2m7YL3CgIgx3X9pOVtTm5sPsdvxMr7mKWNkQ1IHedjIKzi/kAseN1
XuQicsWRf92AZ2TtdBLtK86N0RnQYlfvtZNdCWLrAGZ0B1p5/kBPUvk07IX8pv86BUpzDDrZOVQz
RGj0Q8nwC9TdvRCeqekC3Nue5FZYgozhY5p4Wqymy7uxoKeZAsOHI67GPQfjpbtt4Sad6MQeYy1T
AJLqFccsfYDZQPxlxWGErmd9NZuW7UX4vjy059xc9iWel3O59y2MBJyn9NRWjyHT191m/6ycF9Xg
041mqusZa0kd/1okfsF6bOg+BvLua0HzpTqAhqCGMC79yzsPotGFg/4sYXXJEasvcmb68Di9+CTG
7vVUHd+jJQB/tsn+DPAaPHMOs/oYFBjhoc4uVIauHMpc7QzTWn1+F2OL5B8gPzRDdmgJbOLjLXEF
V8eXGO9kmxo2o6elV2BgWh1DVcVxy7NpluOJ4tuSB1Fh+lKuRaMBspZHIa1SIuyPcCQHKBngtoCn
mx+rj4I2eddrRlcRAnR3iQvzmDskAaJ5qpqZ/nWRDqLaKG0SgzJUwzt319rvxOBpCfG877uCdyAY
039ZujE4NJejvpF3sJqjGxTTWYi7ODWRgzBjNY25wTXHVdkj/CXHiUjNSnoopW69PIDqL0k8LEMW
FIX6wXGPtv/xele3pcou2btBjRgGwibfTqayDWZiF8bhauy/aWzjvgFdmr6GmmOI/P/OfPw4xGP8
ZHJ16K05+oW2GEsYcsnPFnM4j5jfjdLmBw475EaizXNUF9XM1d/qUUYFkhraiZ+wbDSBniezHMvD
oZgUCWTF1oCeLZf7Fewm84z8Tn6kBZzpu6vRCwPupPP/4F4GtqotxIytzEBCNwwSFIdbrttNi261
8Wg1sSckaRO67cmF0ZXR4XAsMtaWcY3WzG7amKiky/Zd3JfOPRZb2JqNyW2FG23bp/3v6FwbLJlm
60qT7AR1cQP7sV5z5ASfxXR3YCLN3Cb/XRzACd2trB+On+UI2M+MQxk4dO1RgdVPj+kYUH/E1btt
eO03KWALeTm1PH+ii8C46Mk/jyOHPd9e0knBzLzw87PmjXCeEqNjPG9peUolbmz5wPjLGmRscn8L
jY8Irt8XQfBusKdlL73I1rk/ioF5fFGcoXBXKG1KYummvvYuBhgKjwpA2VqxWhs2acQjz/iFfRDr
oboNDDPqrAduYeA2B2FGp1KHHRz+BfjEe0pycI6uRHJj6R/g5PU5ojo+gvxVjDWSX+UK0wvW0BKT
yVaNNydAUWBI+f6Lq3+WWdqU0bW7R6iLXlLpGZUBeqcptuQcjJvwcjReE7Phn2+X9IjZsDLnTB8x
Zok1qZgljDX0ZKdXuK3ydyng6YsdzQaDRJ8XRY98aIejjWOI7OQRXj3O9/XaYCC4oEov4RlZhTc8
TN7HyQnabEfhf4lIYpqXwe+I6cdIDHZ/19tLY2pVsFC8Oesk134COgd18WV90es0BA+c7Sg/gOEo
/PsC/Kdjxb8wQ4EoySu1vo87/42K/tn51RuNqUz3CBqofd3BhcxmJJrE7Ul6Ng6VGarWrKi3rxrr
YbE09lUnkc/I9NLssju4JCvT5TlIjC8yuhOR7pmBLGkoAgV+5Iq4lR3knklgBz+p0zQM/PNqQods
zEymsv9yAcigDmZwTq5Q8cGs6j0WnyBkbCQede5Kl6nz7fpKM0GK2fFK+YebqpAWimHfYnsL0O2u
efyLWP+OgWhe19a0yqXjOtVaQTKmwgjYW9FUE5MwbuHBqLQUa1D3UuNwmZJ+RI7r0fRssvPElGkK
Pmq5ICK3p6Gn2kRYMWY5MOfCXm8TTWIsyRh6tlaDTfMWtZPQoVShIQ2lyxHXVUQL1JPMHDaxXbbG
+WbSHJobMl2R6hn7QB6uLCRXQrv7feYOOKtmyRSSWwuaenZ1rLx2cruICX+c6ms82lyIORZab53j
9VFPnaZS5O4r7xP97B9JfZsQoSFhdsPPz7t/TDdmURufYh9IeddvO8pvI3+ejwA+IdQsueWphALf
ok5MnQKZKbhZlR+Qmvkl41oc6xb9+Psoci3sGbTVdgN+RSsJb8qhq64TQXocmw8XHyA7pMtABuZO
4zuKptuD1JFJQk0aY2k9+O0fdykh+mR27dPUqZmHuP0bxJgcGTxZ7wTsC8XgY4QUOHoj0KFxF+LX
Nh//OxF3L9xR7dcJdcZBjMkQ4pvrGqbFADBExGVTVn5gAkQMGRl3C57f70AySpYJT2z0lldyBSpV
0Wf8Xc2e376mL40spdmJYDZvTX7imbz9MBd8Pr6/0IZ2FMmwzNeisXhm2IWwAYMk249QBoo6blFB
LRNdtrWFnjtzgpYbFB45PXK7+CiAr4ksnCWxQWGV879nD1P/GDhSPd4QseiCyL2Y2IHTZjM8W8RJ
tScT47i1q92uaveiTrALTZWseQB2z3xbJ3GXyMsQQ8qqk2e5xNgQ+89mu9aRs+WO9BDZl8hxgcY+
g3vhlHgn22pDxW5nEYk9XrdZED1gG4Xk9WgmMKDf+Aph+BpAuRAI6oxSRwLJBPu+su6e28k5o4XI
ifwEe5fnFKFnovFirxIrB3nhGXPUHCLHj8x3Q+f5QwicqzHKOmOV1XIiwPXmRJDPwZ0Wb8GHSVYq
f4tqLTMQ2ZRKy+9DKEh/yMHw5tm6VmZGUrOoGwv62Qjuuo/IL3uuIj/YUMj9g9YtvtliYju6mAL5
Wj5p9YXqQXSAzV/YQUS9SCLU7Q6vPqE4jWFPxT0PuwZso2rp2nwfYodxPkIAWeeFLONQGFFO757h
VV7SqFtMlt45pDjQdcaHqlXJWNGwJd4uD3i+OordYQHHxvrmniCnFlF/ZyTCkntei/AtiL6oT97p
tyUom0iC21wIEdrcrIH6iggbhmb4ljDosxRbyV5WA/W6LXLRsjiHijkS3dl8VnH8nAUIvWagPPAN
We3xB9re8oLydMZOHrqLHXYasvMt4UNtzhbdfm5C4S4RTkagpmGb/UaszMTK1upuNBBFhfXwMFae
Hn8qnjj0x2wuWHF9MeDqVbjyC0/cOxu1FNnzN1KnIOgdcE5HNAe82MHLn/4PWt2PlI2sMIdHhVCt
TLI/KZVf8N3wCU8RVi+Dd9MAkNcAa2pcArmKTTsZ6ySY6hUSvy0AdNjPDFz6esxV2spMlkeC502B
LoQWhdCl958GDPA640RhL1f1DMGs4LV/PpdkUh1s6+mmPuDbsZXTPqQe53nGEmMJE0Xp03NVfWHf
iaravQ+g69zTsqCKe2NToHi/okEMy3IE16OEQ4qSZVv7JFHvSej6eFsdi127FZ0ZlDPtrsm8bRUW
Ap7yClduVCehzqfVhFW0zOi+LlZGGiUS/9DwhCuMkZfvZHalyWvKWn4/yZ6mavAfHFqTD1XYohNK
/6nLQA7MA+6/VTEdhyuKPqkbdrV0dRITt5XbO1B9ysdE4uPXAGvZZN6SS7rN1nD8ilECnuG0uT1I
xs5MiLtCvxM8f7TbW7kGjWGe8TfW5E0WyOys98NLUxAN2X0Oax8UodzQdEG2O5hPHu67paWej3hu
ypnN+FriCMCPvmagF3HFS8xGDcqbyMzVEHT63qsMDwTPGj7pMCE3EgAVyrIZzeNCeznIqKsfdIbm
hNJ39NuWbOGDPFOqAkbTX6aITwIAEG5JBn5yS+wOnBTC18z8l3f40EkDHPAYLESPagClUo+jRthW
JFFKFimyJqMECUiQbFGh9ITGRME1UE6SNzL50NmML7CZ1ZQ4+6s2ywOobILY6m50R9HXbidlX7VB
RkFNhHajo33Et3+hZ7IEo6mqpYnndX1EFbKfk9VIMhEAqzcAsm7CmOdsRq3uGyN6XIApGSrLBie7
1QTWlhNBs1TlSEFFsA3pVXldn1kvQJQNGHGI8IkdOsNa6mL5tFwgAFtTZye0ju8V5sCh0o418V4c
dpoN7fatrONRhHL8SEin7XmqtdDNwJuE1yxEbEgpVJ+0DfC//5DRqbSvPGF6fyclHgxjQ1p/qmJX
GOCHs7U/wggGKTCoAxa60SMIXKNQHPGMNBoD+cT2Z434fvJXCGvEuK3Pa3u7rSbRCG8yu0WYPpUz
VHDqqTKdRbDt5LO4FlcuiMFSURK+DMqkC1HjspzYGp6WOGtcNwncIiQOx3eQ70oxMsHfKNHv3SYy
kB/DpmJcUw9W4oG8TKdpjm8eYnqvn20uDagqt1eGWoVBBHW8lg2nowRdOJwVu5acbo9RZbh21fHH
LDxoiwZmBNxN/X3uXPnERQt4dCG139NFzi3CX28yzocAGQWyOj0x7ZSBiV4kk8jBAIdh1isK9/TW
M7qJEayGBttxi/RU7dQw2lU11f+TpXanEm3Mi+EZJTnTFORMHj4WgWDGoOyWwRcF7pNr4KuXriqr
e0TtNgkqP/zqUvTOAyL8+ouCKQS7svBscdobCghnwtYtL2KUF2GSSqyMkeyv7XPTa9cn0ZWIDekF
58cJ/QDVJzIwknkost0WsyyGlry7aom2nedfkdoXmM/uuXLTGXAd14rqPMB2HOrlbw5y2EvFTwxC
ioitcVQWpsXfJKeNxqAqmiqjJ1nyWKay++4I0g6mJkbEzCdPvceYHdK2FZxHH7eH7hfLLzbNmsrW
YthuhyBlLatrtOBZIDa0adG3hQSp+KSihD1F9Ur9MxFlfgkGD0sdatVPE8myHltWV3qV8lZwbMSP
FNQU5Vr2p/6Wal2KvzvfikBhuO3Kqw1ip2KIY0fJ/xJHeN3Kw8HBpoiwakC++w/exDwN/fVUCfix
6EcA6xt3h6sDC4kuyEOtMzOP6+l2Lu+ooHTAEQyYOgGz5lhe86J5VgCVSSUZCHagPTSXHQ5HCYi4
1j8iC3ODwQSqwJ6Ee9vE2uPy9pbJg5TOx7mgIvOinv5d4Wrmw2CWyQwuVfjneDHxoEY6OX/4XAlG
iMVyLK64JPwRah206mVNck4VY98oPqO1tEuQFuEglLHs0QduDwKw9lt4wslqzVuvKnOkGWnw4Y0a
+3cSaMbg45xgYCENGpMhtwgixa22g+4OFXVvUMRyq51HLzNkJsuHVJO3ZqffR60lOAmYMfIqu5dP
Pra+RaLE9d4B3gx2/4vcwFtSmERiumYCeKfFrZmA65RVV82vmTWD4tWiAGV85MoyOJFInh9Ps0c5
zdBjBDepztCqK+1NHcLmkAqASEx1mXJ8RCmib3lKX3suXcbGit0x1ABhVD/sWEeDzIqdmDnYUMoV
/PyQ7m0flADGhlk5qSCN3p7yFOHOH3HyW84ShbP7PbMIcniR4NiC0uuSjQZfNxvTUpaYKzzxPqF3
AI36EDmivEUelxEsfXss9Zn9Qh0EbmJjZtkO9KGfTXs9sGX01m4kHa3ocP4v0YgkV5vPQ+EirpJW
7HwQB4ulGncjq0hFSsThbD1+//QAzTGqpEpq7EWhpdIDZza2Fcb0ry6cyNfaXxJCvXL90KzyxKFu
M/cKmpRFLRIeKjlHxuXimY1l6MXm4Ygctg3hiH/Xd78q2kRpXYbgMSeFl0kcKc+coh0hfm1l61wn
J3qSiViRC+whTuer8S1Gwur/pL+1+/EIIpfsOnO0poBZ/vrE1Rmx77uQsCidfCovXVfESW+C5Ff4
ETcpAobWybSbXrYBnWWXdAmpbeFpSpittj5ydEoV/yLt1fJ+0T8ifGeH8ifM4dr21V5wNDnCll7h
zsYO0nJx51yJYHmWFCd/B2PRT4W9/zURDWDXgbODLa8deMdlXOg2mqqGQdwzfDV8rPDKcraOwRbq
1pn4pFUhg1UeRKa4omwuhuWeCxRDxzfR+xFmHqZTDRplutvjyfAkLmq7eZEvUy0JuUTdCnu8oMsB
TKuefymuxcoXmfeI+mGJV8zTdSbcvykRteG9qDrgWD1N6uFLGBncugZzhxoaRXtpqFof8C0H4arx
JwjcshxJjEZB5W+aMaexEKiz7o/NwIo7G2G/U3/P42D5T0tyXb+qRWq96hHFKDrPXW0nOekZGNww
A+pFbuWofclMMOMKKu9FlUZ1TaA3oupKnUmZPhSUwnfbxy4f/3EZITgjjvyKLBBA1bU0fGQHoyDq
efsnvPX1cg3HQg+PTJMuByRDA9scvoeG9nTn4LVet9wDCa4jd+XngmKqXRCNRzphl16PrdBTeprP
u4KSYohv3b3DS633gFZHRT3UKFWAVmLsy+BHHvWV3HWjrnt7PbkCR0k4ZQ0hZGDwde7rgm9qIOne
gIq6uV9rUE+xBO4R2Eznr85DmOQKM+L1PlkUUeikE3uVlkgkxEU6Ux1xI5E7/RM4sDpz82V1Od2Q
KgcT5urmf27tOhZ0HxWVY84lxKZw3aejUCRBwsVukq0yawzGa+8ZxG7SWZ0w0BZ33MtuvHkXnMvp
hyHXTl+4ZtfcBgNWzF8gFUCguUxb6F0aJPsu5pZ9mwfX5R5qkg46P/3Lmh45Zpx1opdAltOqFHCn
aTOAReuoAmHfzP202whmC8FGSEgrBKdHgLCe0g/BcEGpjkXlVY6yccfkfgr0LyRvtxbc5ROFAFj5
yj1am1dHGSh5yecIR0UodR7/fUR0ucEvnyc8sIxgNhU4ihLhlRaWjcQTM5CM8p0L9nAgOmgaq0Ov
KRLOb1Rl7wqbQgH+eSn6bI+L30U3iDla8oPobsW3PjlGukbJSoZW7kajsne1dkE33htr4DEfuMpF
wGPzIFP8PGy9xyDIHihsARNAPQ9o+wr8H4UzBnRAYUzvQYDEIENQmRVKEKvd5bZ0XWTvgZNmSHDl
Eigpx5ty7R9IwdnCwC3iDnwgaFuAxjY5DZHR+gXFdE962isdV71CJFYY7ic/5BgStveEaHQv8A+J
ZZb8upAUNQc818knRu1n5yXCfue9PPMQPrNYEbfEilSIjkoLaLs6MYbkcqxy9HrGv50Gs81hamS8
ruGHMG52zQAOcAZjlqNl8tdMye4XjAke7f23TkrF4BURpnF0h/QEqvaJ3xPDLpSt82CJhDfv/B5Z
AhtzJXpbO+cTFZaXR8PcEyVqO8qDNJjHd/qa2I7iVKOH9VAkjtlBwLhLjFOli7aRToMU7whQ/MMo
yOxigsjZUD2jT/Shqvzj3LMtcNVqpIUQkGuUpY8kzXrxA3yyP/P2xccPKj9xxFyI4FPiuIwn10HR
MtQNFDfUFVdZT/o/zP5LH5V8BywlADlFho2IlJW7E3IwVQH64jR5Wj9LPVGSeLki7rucsmqwIC3I
QXntud4FTsNPu7uGUTIzixvpYn3Ilnlb5EKJluuuKYmkFJlR2UBpd6fcngveUEGePrOfea1kKYdo
WeQkqhr0REIlf00btZ+QEcefA6nDK0dPi5GB1ha56dUkVmtmcIuDGU4auMWdCmhr/GInDrFAq7Yj
SVogXfbhi8FedsXIAC2P6T6/zGyPd3iRMkCK14DNump2C+SMXIyGIhVB51doSiPkHzqYlnOmGb7q
AnsIoAfwkC+swt7ZjQEDUGJuZCBxBnItYkocIhCwgvJhvmB9kN2ciCALbqzkz4GhdayOFVdVFe6s
frHaOpUHL6lg+V5DIti+iiQEL2+3J//s+bXq0VONxIvBNYXC7JvHzgbS0OK9JDf9/CnXEHUaFYny
vNFRuuglxP31AJTsQtk0jx9+38l8r314/DiDca6Dw3mEu3gXnqb6+jhkCBSpYzy0Xlm9M/LvyDqP
xjtk4wBsa2sQyAKIdRk3vUNAZu+ZiLKRDmaLqPLmDxxzUjFjPHNeTdBo4HlmDOJ9GXeKZO/V7YCl
Cs9KVlp+x8u97Y1G7F9PofA//UgNMDtKfLTmncuZQoQSJypL6WKThlU/UKMzKhHAshes6eUJDoHt
bEThuS2qXrYePqhGTiVqbj8tkKgMTZBl+4+YgGofPPVohkRcWn2n6t4nKJBPq6JRSyY49oi2NTmC
O2F07MI6FgSG+VpoZJFSLCsazRzGk9SZlgsIxFElqGed4UiUgLK42yhPHVfAkhLm2MGs+9zRuQT6
zZDgf7TW9mbYKKUDR1Z1yqKhmbGEClzdGct6o8gFfQbFuzM0xDa6eCWMGO44KPVvMS09IkOcI68q
qzODi/SAwSBj6gDq2KtivyboIG+lle/UhcK4RtC9/pZfmJ+LwerJX91FKSGg6GLJVg8CWz40mbPR
3fo8/YYJtse7VggYlJ8Vo9rLK5tgbqJ6/JX9IBeIefcVN5gMR+u0tXUHWw9bmTk1lGv/VfM92NvS
fsk8x0L1fkC7/OKry1b7CB2cbIVFYp8QtpHJS/+18JCJK1D6kXTLFMr07daAiSAK8XXWSCWkXC6d
RPUGoCrdrqj6O/tC7JA9nIs6jCB9M/3+z0mINZhryAYMyCgYdwbljc9ReYLQ/jCqUeJJqLiPVSSE
IINpcGRmM9UnQxhiKcLNjpdeoYvgydQ/v574CuaETzadCe7qxuI6OoDiiaB87Hi283gIpl5YML3Y
9pjjKRYBmJ4qf7UPcNIjey91H7VdkB2oVtkZ50V16k8wYLAtq9z+U75FuxgQUn8cq9wMsVwwkmB5
ReC+k7Med8icIqogLnbSfqPeggtQGBLbdVwX/goQQghePN238JEcumMf6OCw2+tKRrKuV5iM2S1V
WJcgs05HqmzncodaShfQwebDB8EEW+kLbCTxRMjvk12Ac9egY0m1n0QoG4T8KPty9amxpIbwkdbr
s/3Z3MzFmOZ4duUK0I/bOjsUrYqUBunw7JWozqVP17ZqpEAT9QzX8j8O8vUSLgz5k+PsUZtIA4VZ
Es/dhSQ8+UE/ihb77nFVLaAR6BwBFA6iOwnSqWHFP38BDX30n4+igW6Cc+d1rMHrFp/8aohg6pQx
50RP1giAUG/K0tFKrSmDPjeX/B4Lv5qhIb2oSoytNreNdjuuM5+lOJHnirzlKQVdCCJoRMgj1sXM
+LtT9esRNKswc1cV0lnh93u+EFNGU/bK4/LY4iKo5A5mwpfUpcdsA/QZwFjTWMLHZ89TMzfmgbQH
+97rw4w33SG3iwnvSwHSqsRUZPTYsDNqtD49RLDA9EFFwuEL2bJQrPqfof45Rhzm3LP2GWC7hCq6
4xhmXrfmFY9A+L8egxz5nkUkcy5Hf6NUTY6wuol3W6WYZ2i6kZW9L/p0MA7BoPE/7WmG/xCspjR5
Fb8DyfJYaIUAx6Lj/rgvVaOc/049zVk2jSvFRpdfvfQ8KTqz82yD9m8Dy0orfx0Bi53jBwx+s7T8
UfcA4HTT/rgWSekWUmac7qsQKeK/YL4K3RWM9TbI5NPfEK+vub8xGm83UdB72T35p4Ul600DUhQw
Tj6Cm0W78+QnsQh5AlHLNh8dKShvy8LfpXxaocqZU2WIV5xgQI91wyB5/6IEbGVcBb4IhdyzT0jW
IJ94iVUznXzlNxd9Z0PD261m48BURiyH0O6E1SSCBVl8DRDoClCu+Jr3HXjniSBvUBfqRsa2hgve
CtyCHwEbW8AO0JGTWwspPCPHHf+gcYF5grCD3yBLNLgwdlTK52OT1p7636olUMJJQZxRDqZbiIxM
kV0dECsOfcgr/jWf2r5tROO6M7f78m5/Qrd+w7c4cGrdljA8i0Jl1U64NXXTnNTpkuwwFdusGcnW
JXMnl71/BkxQNxBDh7EMYwe909eOvK/Owmm4SamMqNgRHeMcrLKG3kHrmdFNOynHQsxS72HleDvH
bpcGL3xzAzXTZ/hSkGXventlGky3PCg1d/k12gAW1KygThiIBhlGEJmYvfSzrI6u2Im14UlA/Ksu
TKnBannx/FA9IEBejTmYKjiaBErlpI9I0LcIFq0mtycFjEYIjJf3F0duJ+TojAtQuWonez1FdFHb
DKOzWlO12CQrMRkqSt3Z7PdTc0Ow0/GR8pFD/AEa/diSSza6PYAhq9skRM46pwcamEv/Xz3AyXlf
nEy8nR/0yobuIPBO185ieLGxNZplBUwiLJLZx5cQcdjGwcfR/Qn+YhtOkNnMBdO9DMkWDeoMxqC2
Qx9/h1JRtdTl2K/8aRcJTlRTc8UjSzaI2tS9WKcZ31jCTzIuiMEoQ+TT0B4IMvJmOH/g0yNZ6N6p
z4bsNXIjnd6MFYAza/Rve18szo9DyCe1aIBdSnjN6kbNWkTPu9Z323Y/tPEuB7S+ZAZb3Bawh9xT
9AzNBXXjFQ//14iC/+BFSrfUeuJQSgBwTEfFOlCBuYw9+nhBiJkRphCAVUyJvi1sGHIFfIQRdF6Q
kouE5jeMLD4EQ9+IeoGwQcgtDVXVoxldrfDi8Uk8Tc6CxYhFjDjKiVSxBmsvEuPK5haZKpHmE+LF
e1U6BGbV9MwQYwJmx6VtmAYPFeSnki36/ZtFyR3u6APGecn2ePJDKj9Tedk5jWxH9NdLVvFq30QI
AQs1v/GRcsFjfB+XAdkZLNX8em+OeTzEBumcihLx/5g70HLg6aw9UPi/yVb6Rj3iGPoOJu2zqrNf
1P/wsWxDtZJBrDdfjhy5C3yyJ/0LNLFusFzI1SQyjqnb82NXIUlZzl+k8IyhXdUrWQjqCLNMHx0H
lCRAX9T1Tenmo0NIgcof1B5AqhzYvB38OA4fvuuP8bLp9fjJLAVaYWqlhEWbMFnXTL2MHBOrnY6p
DgwnW9+pbRawka6IUmVFImP1R4//zQTrQXNeSzEM+WNPxkZGX4oJZJQSUtyjeDL3d53KoUb51hYX
E3Sfqd26VyzrESq28a1vqTEsdq1fCGP+YNHFNEZwEfgSRx9ibBwBZJvQNidy3mGxsFWicnr+OrL9
Wh4qzJdz2Zfi7G5O3SbVdXZ1PkUlv29GpdUjFrciFjo+Hrb8zolGTkJb2DXSHdp+AGvVfzpI0EIY
oqRVDensP3GwP1vkzcTJpYTpRzLVApMKCEquwIUroGsGvTZlvtNrWFbc0X4nwAPQEZSBr6OID8Ot
PCzqN2Na9VDOjmEQWFZvouzQoJivZoBAHtBqTU/eeJLltnxBu8RFIunl8dthFrD2kMStvxbir1Lk
dMOGUujAOIZa0dARhXaly0B25jsqiC9uhxeUBe3IUMi351ZE4IEpqN+loDQtskzLwn3hYCmlufwH
444aYxZS6NjVOfGw2f3W2En71RvdyB3yLP0Wt5tOwMBGKK1Dsk/gSJg/bIrO+puCCxgH4zf+vxYB
U2uUWveKGT5GDEgI3gkU3cmBgbxdb8HfvexRS4Kgjf5K/ZNPVH9tH1jhxcWe1sua8omuI8Fhx7Aj
OWsKaSohQpdq8/AnXxdYvbQWQBjXclJ6wjA4QTdKxWjGlZZX0mma8ZsOZomxS5iWIhukoxZ6lKES
x1UcNqJxX+0q5TLj9hHGNv/ZIq+VogpWfGCK6WS2t69nkBoy1vmF2cJ0B16yO/miMXL9fHFl+1mB
845HzDT9Rs7K1QXXhnMnyUmXp+2jPPfySGXLi5RORE6JVePEOkH1WDVNi6PRxIGE8DTyCR1Wk5yR
q31Un0Vh1HEaWDDVXPe6lwwMMnDQe9utjDRSY3IHHBGKP+EmPREVMYxR+bFXE0zUXp9JjHf0m6eL
Y8I2BIGi5YjjwFMixaOi6CRsdP/3YjGbKiZ7otH8YXsihRVBqh6KP5sM4ivziyJ02iZHnj3QS211
INVyh6JqHN1dpPQX2C0LR0saekVnaoDg4ahpVEKnxuOUEUNEi/jm0GAaqUd04DgmLreTzid6hpqy
d8u0ovGwmZR4PESBO1ZmCTSwmc0zlOzo1RnGXxtaYgY9Xns/ptt1i/UPQNPfLgUVVr/No4GhFaUJ
f8mAiqaCBgb8xSpXIeEv4QpbMLYlwGUAVfdj8l041S2pWVXr5rTi+MARc+itp4VxCqYcGDwi/Ce/
+udSuQz29mVG024CCCv6JMRV1ab8MayYTN9WZW6gbevKXHEwe1kSd0Wb9twnBq4rlqC74VW+3i0F
NOOTyNwJS9QisF966olmZjy+Nk6eVfL3oOVYCrHr4kfi21J8SPodM9uMMYUlgmraACnFCX1rvNNY
6pa15n+xczI4ZuC4puhArBfR/h0sMz7k6qbr7PMzTd57UkuGQ8ZA9hbdgSpTSN66R95icklc0OLu
Jumz5UHoSxCisZGYTv41fKS6B+uPlNzGxwqwXd1cZ1km/qPzrYzH88wu99HS4JmdckP9G5hvpfcI
uxlSEAj4jIDnjbPJIwvXLQbWqTCxhLCZ9NUM1mRN75++NAO2NtILGJNpdikFi9hGFl4ZzN9Rdoah
Igkp5U8ga3evkTM62k7dMOiSjFxSPRBO4aMlaAYN7QBivSFsiVtNBjFYIvq5qg7y/Z3y9m78H1Gd
HGFbeWz8/T7iwBfirvgv2/XlYTfyhlyuluBbrdVVM3p9WxwC1wnTE9I6K+7uKrRDDiS+li9OGWst
R69nIYps+uQdv8TQ9Jzp8I9HjRMI5YU2yP3sOR5L3czQ+Fvab6xAd3EwDMUjule9bxAY0S5CP/+0
iqNnJqfFdBT6H1tZq8eevdJ4pl0bsvUxZ9Y4ambl/bNg26v81PSPlrIWEpy1ovRsI3L2U7Ac8/N3
kfyNBQtlCRljugP5uydsJWdT27ha5xkT/KJDNMIhq7R5p4Mfo0WV9qa4FqGs2yXyoR/BF8MhYrTk
uFa1sKmyQSjH9orHcCESan9J2huT+xsYuh3URLhYWxuMFsDvJm9o8/aH0FoWtlJjI79S4qnPmTDV
K3WE2UcJlwyVXlDYO9OqjMar75Dx8N+m9JlXMyRypB/OP4NXFBf2Bdkh2dLOqkZNYx5jel9hnLfv
iYDAWBSpKv2ZU4Nrq/h/2KKcUrF7pJmOD6W+dmbXtng7nrETRCo8qnsrMN3EC1NgeriE8NfEWOJV
gLAgJgxdjQGVyMsL7eEpq9XSISiwvuzhd+RtHzfAmhhx+iccFP7V5vRUT1Y9P3l6noHV9mjMxmsl
pE5CP6JvaVM2alh72mrk6s7ZBjuZqz5PyKyT8z7Nm+AtRjedXba2wBOIntmFBNIuH7QHVO2SMyxL
/GFW+VYeOHBZZsME/YkLKOlVYFu6Tg0XfPAZkYVrA9K5z+DHw9krgfjeE7SKDjjqDMbzUGSUi5BN
9cFQ8YYluXREuOpJic+md1yg+nYHqWTYh7jtKhuo1/UhCxx6f+7cPwhy5J2lfbsCfgR3A02t2FJC
pE93trxLAvA7wlB+a61IO59sN5Ujs1osr0/aAgADGTwb+LEFgikJL92nDzGUitJ7tVkH2bDQ2bai
+KcdbDM/zuQ5Mm+8GZE+ywInp/eRFkDCxMDM5gesBDEyD5/l0DSj+q2vPGxFvyEJ722avCuadcRJ
vhr6L0B1/4OGfbpRS8jp7J87UcpRVRdIsS5C7oHZAQ5suGMEWrPI2Yc2tAh96D/NZV4PjM1KFaJm
N1mTEcH7gZcPd+I6C2Gzn6P+IcnlLlfIa45v1IHA6R7l2fxXDcR2UxzcdW7VbbITWBQF93yyLT/J
uqhO0+qQ8usIFAVPLtYYHddsbCSa0hAp59Oc/jnxPPEQP1DWdP65xINR3WuZv+7q4AWvXVcv2oWb
wADELzCCXd4TEOKnt5Z06b9GFG9+f3gbG0PgU6iK9ma4nNwrIGgQGyPIVOHihpmu6ZG7mOU+saZg
h8+N+N/qwHrfumF7egyBXLcPNgx9CsLHWzh5BE8NbCk6xnmwE5mTIrHPisufNeAdrG6ceE+uy6CF
ySceN/xzoha4kiEArH1hGkK4QtpKmJ+HFu9bjQ86W/dhGFBNeaGtL5pY6WP4GN9NuLi7kNieyynf
2VyHuzSOeRnz6AEt9QY0vFGkIRztVbxh9uDGTse1oOcF1Pyn0JECazjpF9yZLhky6xTRLg2Cf1cf
HJU2DQgs2TPTJUBB7yuoHz+0VHTs8eQmClwqTnRLNU0S+5sd+2diTAeYSi5kLGxwSPefdTCBkb3L
vqoD+QBWztMvwfd02ROyQZ4Sd1uti4XnGf46Haf+OeelTp8gAA6OlPVHTDKUVNZEodxh0AsIySXU
JX/PEvlKa0DVfBNU+W7UMV9TMOgWVKUxpgwQPwOJtpak2ljzzmnDA0YcZdRfAX0KG0MTYkRmMsqA
7M0X6jvnebDEz4Io3aDvPnzqiISEUhU0Hw5i4oawWkONj4gi5ut9iYAhnJYtXDToUW08543WDutR
yH+DqxpDGY7bqgOh8oizGmeQnUMmyXrPNQKfNgmeo7HIY2NHUysBFq8iT2BqK6RUSbtXagjvvRUm
q5qV22yLqKo9+yHg/wr4moHi+IhLi1HTPy8GdTrnaUswNiqmKrdlxzbrtDIR7tlpKi9dvpcqggDu
+jOxejVR9jlJy7DLyzfN2rCY4DbJ/725sPYklXlidWTLlAaf8N0k316RMpqFfjgV+afBzmqh347H
N8sJIRyRJwsDvZpTD6DyoKUgVzKxIaTZ3aHM6WBlImcnl5ndgMSnJjcKq27isFA9dBJxSxdjmyO7
feThiSC7Pf9CMCJd1qwk+3gSJLZy2Zs0n/BsNuEWYGzfrpKsHOnvmqS954scdqCQnEMVIrUS7H5C
x6uquDrLm1amSENkfcSz55D1+b0cf3wNfEM66Nb9ym19CKvh9El7hb3uZY9DDd+5wSgECTQIpdP0
XEPPgt4e5quV0KNpA3gAG3n7fVmSPOatoRFXrhLWek/8sxTtoOuvLoiQ28UO6Rcl1OnML0+WJdH/
yawM3cEEmERJZzwu/R1LP/1apw841eqpiCLje58qgYIzvYAHKhp3kQfImnuhzd3Wr6hiq0paYc4h
09s6jOVWjtIwSA3fSsLRKlbqm11NwnniKnRXWiSPJINiPpFzkhS48Aj5lyE14Y5swm7LHwUAEmZb
9KccuOFLix5A3e79Vhzh96XT6QJHOuOGIy2RSsf1jEtLS8t9PRng/bGdb9I0GhiL8pTP4qzD06xo
jPfcWIQxxOXjB01rVm9B2mUN/KbM20VnWnb9ZxiA8rynLd0p3RYbMDgITakkwdjMjgOpcEF81RIT
U9Dq3roFFk4UViKstPbjE9yMo2TPq+PNruyV1NwOdv7vZtntG3agqSMBnh4LXyse4wAlsx3PJHIu
vl7GNC2x0KF7vmwCDqtPIbBBpuy0D6Gc0fWorqB6r/QfCNNinuw9CkfIBjB3DbrbtX/3ofwgEWbj
kbv9jAHvl8hyNtXzH3hj8OEAyb2yj6d3qMTpF1LhgkGrVfHQ+Vka3dd5O9T8T0baUq80TTFRd/hG
dsl+S9YhHek5rhNZNs9d88gFk6gbw54U9do4FWU3mcnpt4Nl4DApFL2MIcLaA5BYLzW5nUOQfLkf
agJpL/Br3DUAHjJdpJghILgefHWPPDo8mPUCvOsjsFo6l3kYZCKNFTdTfmEcjzRiDJ5dmqvTJgJH
KERDqmEfdYt5zXH4R+zeqgocuER5JCPXqNR+tNaX8n7PsV+aP36HN7LNIxG2eXCJZ3uZsG7FR6Ey
5OBsDGUYiNdGqQBTH8WAZSQIFbeIer+IskjUkiTGYHkydJtGqopwG1QoRRw4qqsV/U2wSjRVG0MU
QMM8SoHvO1ye2K9AkZea4F8OgauYScThoSt/XGN4CQpT8SJpYx/RIRLbRIFCtZCSTeUxYet3nSiY
V/riiE6xR6CPMdxCThYS1CGegcx7EW52zH7Oe17bOQcctaod59WkuXpS4ikAgSq9QvLoezumr44z
Yk/i3yEHRPH4C6XXMHVAoVYj6CBfpC1GTTbXdkpitvDO1TF0VTT5tiP13nb5jLTKVM2LxEQKTZ9L
8BwWSOUMQm/0DRz9U8wAm336aVlOhWhG3nQG2BIwYdQ0IkNdXZQhvg/OyJ1CsKgMpwyukN0UGP2O
TuZFyc3PB7/47J8aQwfDlQB6JupUcHUPDJS4i9WUJUC3uJXA0erR1pRP1B+sk8QgISw1Q1r+ChQS
v4yxwovTPVFqe0PTS1ebaIDJtIEuEl1N7NfZ29vYn5dUM9fi3+Wa46vhWE6ccMbPH6D05AH/5gS9
NUb1nafuiuDyaFfA12AlV0zEfs5rH5TVsjq/JnPrBxyTP3zDj9AUcddIMBSx9eOGSpwszxs9dbom
Nd2W1XIcyByMPza1LCO/RmKJEQ+GbyRnWvH5UnsB5eUqm1Wxo9DP8BAc/jJHVOiQXukzLIXUeI/n
45emPCLrEfraBZjhBib6YVf1oYj0bhhdv00vFw+8YJKomdhQP7oQ/dsvS8aesXZKsUSTz3yitMho
O0+2nwzrLffhFJP2ZREBw48C7XG3firbqnT53UMNW/yF+deVlUb6baOctmdclJXtIUgS0dvkCIcx
uoowHDcupDdua+gr7yxwg1uh+dh4wotQOLOAsugH+Tk790+zFHY4P6TKoFh5AemdeDSYHF25Q1ay
+Ec37lV0+Z9MT3ZOsICidu+bfkKqtf2Br+1yOKe8kzb011KvF0R65/bwXQbYmgZCdKrxooXg7XA1
oCLWlh2cgNqP9jkQxzsFNC2u0+/uSxEAFCx7JqrhrXCUdxyFFWsnV+3jVrkWTK845ZOPGA4G2gi6
/n4AlVa170TCKMVJnCgOMwePSJxmKrlD3lGzzokHW6YUuY0tDYVL75mPTW55M3U9k8vsVkRhluKt
3D7OXiKQ7wkve9WNtWRSjTqdd7VEQDFQzkLu8sqbD6nhFENzCnJRjmWtLmwK62hdTyKohawX/nlR
zJ+h/gvvcfc4pVMSPapkHLj3PeeWhUJiWA1PsfgpmdguMJOPO6No1cCTLT8Op2UwRZo6ptyb51Ir
uui2E877bZZngbZoLfBXqO6cIwuUUVewZmuWJbDPxnOssDBs0+5/nzBGvcMwvAz6Pwt0uLmVGC55
BSx2j5JDqUAc4e72i3EglL6N8oq5N1TSbJL5S6bdaabPG++EbnJAoAX3gIFPI9aTvrmY5xctOV3H
ZwUEBlV6RCbAHq2X1A6lGVhb+UafdMpIeblW4Bzy4Y5BPseaxVL2rgD8bJiaIah4QZU8HH4ANorr
EAxybYsi5f1p4uVo9SALaRubswKtVz6gRoRpfYfwd334r2gxj+pbRaxPTvwk4VsnUQkCsU/7NeBQ
HXO0EbKfkT2jhkxWasG4bRmvhEt5dRujuIxPHUcK9MvHgI9PGXTYHJveYdZ2dZTe1SJs9lku20e6
Y7VRAOQy5jG6b2cLEE4vX9armsh6n+GR6ugbv2FTbqqn3rP6doOLCbWZlxpuNrC+gTRvCc1hyqdk
ZSC28cU1vU96GfH6fwCP1ritTzuOuN/SXP3X5tXdXFinqKUTY+xjIAfhtDGNvOXy+/3YX6GimaBP
Dnw88wsWSeCRjpCgK9tuBf+TsasmGcDuIW+taCdD5pUi5V8T62O5MYskvPVzhUf6s/tGpKyREWIp
BUOHEQqNUHfaKyXt9s5A4WvjnHb2J0lV5NR86E/0ay7hu7i9UbspeRYVq8QpMOWtPlIm8rZXm/8q
PFLiaAdduus6HFe14Ylq0y1ozapyOaZ0nitVyO2YcgxJz2y14DOcqD5k80Ki6ADeqvNiY9gZRYKY
g0O9nPekr7fWfXI/p1iiol5pbhOw9fuS2FMLm3wkb74Mk5dNQe2KGhqhVx4W+uR4h4BfBmv+8TZD
0xZvoZWFnAymYWYOU1xfZXvo7abpX1VtEPq4OflAa1WruO1O/F9EAD90byziX8RgT/cjlplryoBG
t9JLgFa7VLdqp+DkyLNJ/yQy+HFunKJQp74cpumCNNS26A1HIzexkZhV2XEiQWf7dg6dqn4Vj8oi
L9hlx7qXlSWOtnjwCxWOpzqgC4QXf92PWZm1nqTigia26KEjzLmdANLMmvKCUAHIXexL8eGDTfdX
4rrRj+s6Z2EXiWYyOQ1sKOqkDKp9hs7IpFSXUpyBuD+m3yCWd+KHQ4RGyKXm0zqBdpsZHLB2jnoB
n3v4l2lC37lBMI/PJjcS73SaY+uthny8g72LshaJDwY6wA4ti9sLaaulrKwxbrDTt6+7BvUjVbsG
BDbzMqBr9d9NTChVDgQrVNQVAxMUqOMBsN/RQE7hz18jqT5OjZHUXU45zd/+8tHYeJtxcNCho0rK
HwU+FvQI/HG98/IXhjgW1tESqExx+LLMZ5E3275VSYTMQgUqd4IRU+q9aIkbGy3Olc1QyzVcLq6v
dl4qdQMfpRLrsMEjF+VImHGSuLpJc9QicZcRYGOJVoSGjbgnXVt9ieBFKkFkg8q/wp48jlHWYl0E
jR4X08MLsEKM2rXDnyfBDh9wY2jwrV+RlTcQ7G40lPWHxEW4ywuZbUHXbr/dkCJHc1u4d3LPoC/B
qX79toqepu8g7eOdTzmQPJz3zOoY0g4si5muKvGffPRQNhtRaoyyuOcLEFqDngTUM2PcYkQIAXN0
0v6QKdDrxGyFpp+xTUSP661wmLEwGYiT5MpLhY2hUxU5wHgLoisyzJwxg62L1HJP3HMzri1XFe+n
E7k6lZ7uJDkeemt14RLIsFGiatqvhfH3e6tSikKdHJAKko/KmGQ+zSkvv49Qah/sBa6M/cyzwYoL
KxlH+/681MCvsUiTWSNXdGEvZ3zwFPVPa2l2RnUtde7UFsmWc+fl1qCCqoDx90F/RaJDU7LJ0b5B
NnlzBw4tIaSknap82TIl88YcNCCacM4pyfgqNJMLiGnMPKpj8eokWwL2wS3atd7ZBBDr66wMm/Q6
SU6znk2MPrr39X10Sf14pXoYy6ud6owJGVUOW2wQTZtg4ahIxvm5Vdr/Q3VZwMP0AOLUuR5KxpZY
gDKSh/OgG61VSBJGbLNxVCA+7Vna9rHhjSsueKZ86SPaMq2mLdLibVxPPq14Gj1COg7DTGdvSSJX
NI8Twqc4ZiaRPqlL6q+VyCOxe0gA33Dcjj0cRELPeHEL7WuavOsADuBiSDtPe/DZhELz8o9M121N
+PImaFPKIFt7kZpfeJxqqfZ687ji12LNRUNOAGiza/e4rcK3t+xB2s9iWQRlDnZHoIExil+2Dab6
AE2SejQEjXiUGBmDQsyijCrjVdRvv5DyEhrxsEt58zCJ9xzwCXdJGQWexeDexqsE3vAgVcpw9IYF
wmNmCXqAwJ9h/5PPXnE9+zDsHw7OLstYF/lyN8oJCFa3zxHp0rLG4JBebQRg5vBVtlrLYjs61UCn
5TKryVYpo1byKAIXoB4aZ4GAlH3e/lMzRmHFKxLcXNQdmdjTUM56d9P8PD5B3qeDs9mNtoGfhfTP
b/ZXfnLQUFl8BYkjsf0fiCvp+UROrkRzGhajdKFL+2+KcPWngHrWHiBFzLKFPxPZTyOJHfwpbScd
szyOH9bUrwPHrPrsSjNbaM7E9ZhzzwBIWySsOnxf+MRAopVUxofdnBjxn/eGt/St6bVYv4S/Q/1/
TRJ7M2vJCN/lX+eMt16y7gSJ1dzaleERF/0CJfj6E4Ug5NnTHN5QgDcuwwGKqM3pER7SfMtPVreq
3Fv78X54KXhPRCdTDvoqbqfW74f9Cl2sh+X3PmN1aTHDuW7dQHf/va6hWJyo9I60VEVUJPxeMORG
TBZCJhp3RjfeS6lrlTOKyRzyQP4C5kMiLwdqiVczbv7xB60PwEOo1vq14bjeLYjvGK6kdTSKeJoL
UUyvNJM4BDtCJ/KsFseiE1FQtDjsuph2To+3kw96ODoNQyrJWmfIGXMnmyfnvezIZ+j6G9PtTeiJ
BSuWm1yN35Yia0uliSOZS3iaQA0FP9bQxP56J7xbY78QawEjnkjp5JHZt3xjsS6A3+x6o9zCUMe3
GaxUISVGK7v5nANmjUAAq80427vldNzjnK/2ZKBQgsJOKcOcxpVvefOl3BCQT3BjIDy8BRCiLinC
w6+3CYJIW5e49SUvpiY/pzQVBkLDyPG3RGz4UET+pki70Lw5POxx1PbcMla0kWZFgd3DnBxWDpLL
JIFDDu7753gHNQ0FHdYsz/owZTgB+pTQJovqxbuMdQm5ZRiPacStDJXxBROqRjHtLbGQTBf70DCF
r37wwVCakTA3xNMtNRQZ96Eax8JcxhCQy95ybazLk2dwnpxZ4p1LKTyU6ktdw4a+a+p9ejH+aVPo
pHMeKCLDFu6jF2JAymp/dRDSE9LoQ1mZIn90/XlMfUVw7iXGltPQfL9SsmBP0zYW6KlCqJtGHwOY
IDNUnDJSUAgAhj2HIwLgLpZFCJTwcbbQjZDIfFpHGlgsBILNc4d4BkWKU8r1xkCU68uFoCXdlEZZ
3b4Z0CYGMhQLX0hNLNuvBYADPfvFJODdT7UOI9HG7Ms0l5ujwXBBUhSnR6o9O4S07Y+BrQoTscKo
O9OX3JT9z86QB28akWgkN+E18Rxrl4gVRQwwJSc2+RU9NbegXDgRVH7pmzmVIOFkaucG0gkQ1D2+
iD2BMbwNtSX81rOo9ZzFOSfGiNwNONqBSU+0l6Z3ORWmtGl39engoY9jm8sDjgh3gGTK2Z2DTWU/
M04MRcOJWwY2PPfPVWH92mRxtjwYi/fAzusMVKLs2ucS6nVdBJ45otOW8xA8pxN/l6gORp2imN+x
1ZEyba1m/ZLdxDF413EkPfRNp7KtUJ0xnHSJ0h4zZlO0pjRoFaGWf5s1bG9wB1ff/C9rb1tKA7lY
09OezqA5F+c5tnO7Bre/u+79+9EVJVjT/j3i4y23M+sYLhOhbvIzEGFKAttSBL4Bcm6YcsHUlVcf
r1PhCHlyOgeMTO9A2G9Smn3dzL40Ze669LRRGRhXGp/abOMmY0PlEADCke0e0MN1ZXgomBITHphd
VI5X9+1rHQPszfBjLa7Pe/Th2L+QJ3/Aajzt+HLpwjIQFTQ/vDhCijzags5IusykJZsvmex+BYwG
8ez9N+02MByynnojL2zPF+OkEGXoSnWM9dcCjwVMRQYLRAyRvenwg80lNn3cfTeboxEMNHBGEuX8
Ttm2nRtg599JLd8a0Hubl7TMrldZXpCKcjAslMpP5aXRbMtFXryMQry3wxc9FktmxZMtbAC9lIRs
XUkfE1GMI53tlYd9T2n1Go7sXeHVzsSVf7YgldX6Nur9LkYGj4pGseWaS1y+/wyAbB6YMT5EO0d1
yeeD9Sm17jxfImYVbeUa2SuLiOUPBeZKsDfSgKeEaT/5qBJONuQFIkVQsv+E5bxTYqFVp1/VBxrg
4hNAGDvDV+2EJjhkjxI1FJMWO075HUWwl9Yo4JuVQPBwCtCZGdYpIPTs1KV4chjI/ZoUr72EJ/yH
giLCr4QSx134lJtgDQmYOH2H/D3ZZ5NRbQzaKC3wh7Qb99b1cbmdqgjYQSVgftX+cowqshrDawU4
Yq8dsVEqFLHPKRzlLU4RfFYYK4ZGAp+vEHqbCh4OZSKyQuPbTGZ+x4NDGzD7uHnaZPRBIujgUGAl
mItbqv/pzWa7b/IFS9qbr1/Y5weZ9DhZPe4ufaBlK4WuPpqnKGj6lI3uUw75XOd0YRCuWpno5d1p
JvmW01DsuLvNJ7o4pX+c+tTFmAtOU0F/sixb2t/uXfasC2JNWk8f2G48a+3FGzAQz+s7hqCF+Afa
XYZQA7DH/OfpiHCvoDModEk3mX7CyYf+q3RPoSUOfw2PNIP2hdQfJBg0g6G/SpuIQLomFjczUx38
wdX5e1FTVJ6eRG6zqi5fwerlWPBkLqZ/0Opi6SEn46h1lTqZtgYKLoPcOWdN9mIPVCJBexT7M455
+dBQ6KjjSYu9lXI66zHvbV41PBHbqU8RM+ed5ZJywYI3aIr7FJvfE5jVPusMK0DRcQee131h3jBZ
a1gcuvJP0ELlS5LkaTu7NSCF9syKiWCNSPwrddG8DvEaQlARg3g7nLyjPx8r0JCWKLW3VZ8lum05
K/T9567m3jB0Q2ltSVQ//mUz2gMPz0zhExmDmcL07KhdMuBILMMYiyOlgffJUp2MsKpIR8+yyWug
rQdG7xOL4yX0ZLXdOmQdoVNsbl3fPRCjJy6C+A35sfRql3ebbM8b4oT1DdKjui9yTYaOsM3P7IIy
XnkIqpPQZEnifksXBN8AQ/zqRTcBJEmkKM3FCN9Ka6MeCDDqnLzxY6B+FML5uBiUrf/8h7TCbO7v
1iiQQJcQdaOLvUvYaBxm5JJa1csRWDeajVkjimsJ5WoFCkLCm5q5sf+oWI5HOWSrKPLYzwH+C45c
l783h++MDWRmAfpSdxU/POoRivCQOG+e5LvJzbttAgJ4K42ZUMRQyO0s5Hl79f2tyqP0T6CBF1Ni
tkOMtNJXNzzx9sGtVpQxCETJYieZBfz2YSYCRzBy0H0TecByVFQWDEH8XhFYb17fKfDOV/Gj7hUC
RSMvYpN4dZ34i/xVR+ftec0li5HXwXYTp3S0WtLR+93o2FRPNzijdtRBZ8SUPonQQ/re8TGrLFi/
FzMzYOadJTNqqkbDCKSUlZlAhZ5pb0LEEarR5h7Cm7ejNPvl7zgbq0HcdjDbBxHboQ58YXPZlzeM
lw9hSzXn+Fo2freEgLnxy+fvVTfP6Gb6gxxpJsAIsY9+7T3EMgoem98QAwD/8FoLZUwHFHAuM3F7
DSAP6c9rbibtrLiU/q8oqJiM7zjirQD83dNWW6gFS4kucYt57/EaaN9ceGP2dmAzN9ek9vM5y2pq
ciYcTyJRJ+a7WIIEbA0f67pqehc8b+/CqAOAEx1n8qsL6OoZH0PSo3mF6YJYNHLkeS+KQhmXVx9c
gS6ZSX0zkRCncHAf4/eQpl4iqUrwtf9hjwI2/kObtO8Ne9P5jnwEg6mVMo+5gCjdgjtt/BsSEPzX
qXXvV4T43w3kskN9bMftEKbQIIEjNFz9FAuCgLYLDI7F473jpAuHsNrHjriEsaZiuXbFsqBeuXtZ
dNrINIMyF9lOj4cQ/xqYFiFOd/1hEBMAh7MpTlzZGLCMkvMdxOPzt53PK7z+SnsGSdlbHHYEMMYT
e6mt1pnu0DdAgYdc7UXG0p84Us2iMfMYLIY/2htES8/qRo9bmv7xY03gUKU1gne4O6pW8IeCm/pP
jJEEK8Vsx4J4Kgp9NJDA4UrZ9VOTZGI5PNjMjDffRCEuskjb7MML7Q4cV2PguzAzPQSmQM09MQLs
hGSmQ7qIi85Gv96AGagzfYkEYp2xaqjD5tuDQCI6VqrIByLY49YuYijs5dSwb6fArcNWeX+Z8FYT
JUcHpkqWTUQzUBkZNOF2A2Whiift9DrnnLIstQqg5GaXX4EnoeRv1A6nwa7/41G3wS+IyYuQDmcY
sjiP9YEja0u9AkxZ2j/W+C4mSoWBiBIK8T/LMCs2+xZYiADN04ZQ7t2NIll0AKrw0GUQHIY5KdWD
xD/+6qW8Ai0sVcvx2CONVEsbv4AB73sa8g7j4EkhjWK3uamqulVNz27nRGi4bb8fN5XLdSf9eZMJ
v3Ea4JfyZS7FoqX0z8iICLnaPlLJMSLk6w3sqbevHUcZKQyoUGAwt8LzMHnTW371nJeb8ZPDk81r
4cGFh8DkfBv4I5oWD9vlqLixDAou30P6NPIZJCJINCHDLWl5SPLttWfhr5DzS87AS+vG6Ug/LXBo
MoQ3IUz6oL0hizs6geuR6p7Opdn+FknvR7s38XjRYIJ0tTcVhjH8nO5u/EcQTM+pynGa/0B2oz5Q
l6l7fkYtTtcikZTQg1DICf6IJyOXyaAdaWBpbigLqzQe7MEjgu7P96V0BchOpSWqvza+zdWS8XwB
beU1+KugCXQ9JOilAlyVB2I84PvgMQjyDZdgQnwdz+Ks88gzc1QSROo8023jACd7WgGfDAsSrKeP
5i4k7XgD4oni3bD235gHN9QAPfolD4QUd0aFaD6M9j76CQgxFjIvgT45hTdOQPCS76xmYKCkxIyt
gjkd1wyGBH5vjMp5PLQIrWzOrcYiNdRdtVmSmBzY06lCe4gTkR1kxnYznNQHiRwlfE4zkjJyXJsE
UimBrgTdJO+UuDWuPPu/4lSJDmqvahyhosCofI8JYhEYrmwjIOGj1aNl7FQIwBTH7yWmkQAhNNAk
uBTV9i3krpMoyZvfFw+EHfaJLSDsGM6pFdl87EJK1YdRTjR6K7v9Bx3KO9Pzh0nVGIWbzuABURB8
OssTbSDuiVQ7UXl2+ZpmcxoMQx7mm5KTAfmtc8d/TL8DOkO+HLZfwLhPKdDk4hlwK5jjq6QG6zY+
nBNnO8QRL4ksRIlfZL6Hc70qpQdGulc2XbVALmyS7SiBk2q7OWotZKt8FmvUDbUBnwIwMps5tF9C
pVxAnL03NPvTkF4YbusCDhWcXRcIa6YhUbOY26F0+86u/TwowzhkOhpzIxCb/1mxxvxPBl7uSg8q
IUkU5fJkuJl5uQ4xtPET8DlBW8HMsAx4LS1UQlXGOsD72iFy9baC4eFcZKXLS7w9T22Xk9wYoHcK
OggpySCoeIKA6JggtsijhZW1xsT/cnTQHLdYvcchrkpQb4Xc35/SCb2IM/HG52nWFLqHHjXwrGQP
c3ZAGkVPPsmIH97wr8uWAazA5s6xOtxGTG7kzDQvz7XNAn+HQjOYQ70MhdosCSlzrLZKLeGlUXbW
NRjaKSx7erVjDDtoYK64KizFRq8na2kZEU0gtXeV7HZV2mz4CjyWpW1Jd8eqruQLvekJ/WCle58j
ztWhX+nw1coQU7ZDMF84qsDC4fwiaWIwnkiLFD11GpajQ7w3vCHgVzKPCOCol5UYG+iEYaoSEX9u
kVMsKLjURa34HoKDIg3W27cccG10enJAQflCMALqg6cwcitm048CSUC0vPDE2t+eXHP269djZPv6
pO/Jt5YTnjUYp+CLzUDiukHvWtfAmcIq3m7nQR9xdmmsispmyfuVrOX1F15PTpjPK0KljTiu03S+
H6YH8tC9S5QgeIK/IcIwxdn4JZy9OQ6LhutMKA9fL8xtKzbJ94HPyn7gBXIf8Mx7aYnmKp62Wi9/
Z5XOlv2i1rEqqw9LbHyMwwKnXkCj2cN+rq5iX7oRPhyJei2lHXhkg/RINV5CDXOqnDd+NGha8eYi
MZ6c24XgeDansXzxY7f7U3y5LzHqUEPBzMD6HsjAC0vs8m7abQ4SNVz/SFR7kGSZ2M9o8qIwnkeh
KjUeR2RkfPWLLwxuYMub3FvBDn+q+9gopDNsySO4xsQLROPQdQTwDK1K2z7UZPWJ4yf9Yn7Z0l/a
fyGjnJgEkAl5A+xUnjb5aBBFNDdmdijibtp3ArkhVth+Ph8Jhgm5Sc6hQz6ljcd9xIXxkJon3XSE
9vRa1wxSCndMkovVmpkaNFUaPzD83BjlWGnnswGeeKD0NRbaEEjJECtsQm0UA5Y35Tr7ttNiZI5m
Pq3zkmRqMdRXf0cEDgMM/9LZMUTldddSvI3CcWxrMIYdXboYU9Lxxkdlk6mgEvkWSc/KQ4WgSpHJ
3UsakI0lrcmtLRaQVIxLRrwkVEu/tKBFBv6nqVAkAQ0Vb5PnYxG1Th7Bf5xIQJzHNuYqAuuq6UwK
5txXKDjwYqIRlcKGZKd730RFZfjy4BORDWlQn67A8VCoPyQz+0USr4G/d1FS5YSZJtyEYhSObZ2L
iNNkYBeSCxHXIFHzBwAbam1LA3PmBLChRH2tvcQdlnTnUK7LR+SooXntl5H/OxXhMhNYDyhHQTS1
A3nSeRLisPbM/2tSSKiqdhdG8k846a3CV/+oZz75tS4ix5dL8KXZr7vxQq33riiUYH4/Oj0W3tmj
hDBYsMmalVxpV9WjKs1fCYcnQl3OGhWLrvhpTAuGIzIgHYq8AnsVJSO4P0GqnsPU4UzrdaCNIaKi
4sQrD7qp6YjLpWuWMN9YyozAP2ArAxUR0LIH+yH48PEOFQoKniF2r3QnUx0RzQjtLuKzsCjhJP4O
xA6QklFF09S87cYIYplN6OfQvNGq1hjmk+WLUq0cZQtAedR/oC0OiT6XSrk2lBAMlmJ0IEXpJuJz
hwomZkJ2fYS4gycMxUyUKnd4hjNzI276hHtTa2qsDZYxN4Fwj70BPlwyl5zZNEA27ptE3zQghiOA
8uPUrIazLIvPGXBNWs2n/CldH5/8ZAyiyXfMBTXTzIrGcxKesamgXiZ+UW1V/Yxxs2j6hrDmWl4x
fdzprXm5EsLQFEBwm4JBPnoM1UzP/lbMKofpRDSksrFWAONCO+E7xR/uLEU/16j7CCWHhPNdxewy
/myJQOqdx5XZwtSy80vNPGlyG+bB+P6ODfb9HKA8DYQz4dmLCUqHUDB+stT8ueDATSCxyvjhMrfp
IwFtyFCztoiiZMcY4olpPB1DfVHcwjQ5kJ5oIaF6DCvSkDHksMt92K6cH0xDdJaMQev5KXsMDmbj
0TDwWwAv2SVuW1GA7uSjRLFl3sW7nSA+yg/Og5T2AASkrIkhghvG5sTDITJdFDBmYqnGZR4rFjkI
nIeC+obMbFaaM+FJCxjScyxG+Z+FvxK7CytLCyvQBU+mwToGB+HL1GbFf0ScpMU7U91IJysyGGjE
2ct/hy54BQfEZZSWeteoyEfqcHV/c24XF2LzfSwnBW1M382JGN9AoqTTdGIUGLn9DfX4A2Pef0XH
gcCksvw02fRpzIfKBzlvz67OFq4R7G5F+5xlNcYU3/UPuvgbaWk3evrNtmXsqUlXiGwdrgas81Dd
Ms4VHYszRo9oHOrvdGG6CvlktEE19NZ8mxNf2i3aHBltCiCl8HkT+UohA0wJ+cbiQreBmgyZ/ZhE
9bgZfssS1xmKr6a4StYX6B6K0KGB/Z/uR1iEBSH/nPYuShVlFixflaun0BoW7a1TgOiNrN+xbCwV
D0WD56i3ct9tIcFQ0V7Ukm9iBCzenZRGfD73hWKQy+ku9V+wxfG7sezpDnv0aSvQZ8pmV3jJvfYy
JWal3mYrcEgQ6ewgA6qLkOWmFraKNxyoZQ5ICC4DebhEoAITDJ9daV3XQnVumNGunuJD/Vg7ddVp
EZFBP+il5eLftvgqYEsDQqz5Liamse6AmKEUu0u5QfRE3PadM4xzWp6AjIS6M9qKBLye/RlwUwp6
WGd6zAUBvwi7mvnVD5OF9Udel+vH9Be0N5hwUpRJ6jaStJUqKHqyh6ofrvD9xgC7UPDTQKUa3H+e
szfXGlgleahD67QI4uyKft24HfbSPgwEB62YqVs4LuKjehSS1XOG6xk7spYnqGMwn/w2/n7TxfJm
weuh2P8uAOEyvGzrrjPLUPsxV5A1dNbm4orZ5Tyv5mzOwz8C9Q18GH7OU5IAJPD09Jkq/nJBWCoG
8h9Z8NHmzZ1H1ARkT2GQ51+rzKgY6cxM+GGR5adVheM0Ho8biIYAlhton50oySv3hPqFENdzdwUn
mmGouUKi7UIh7+JIWfq5jRVpfjuQLbB58dik5EKpzeQ1p88sczYCvTtxDSVPjswkA59vNaIWPLk4
VXDr8QCX2wdczh87LmjplPmcqQsLKinmAzG5NbYqSl6LNIlWcSpQOPCfXGta0Vk2459ZVeDGN2wS
XJ6JHi2ivXU9CuteTA1L5uTEq8mY/00sHJ9UK4twCQCkxyQJNhbE/6dfD/5SpQFaw1iPbIL5Rwap
SwHpeqqPNKYIQxwZuKk6U09dPmMofdpgKp8FHq+qWXDTgODwukiofVZR0SwVQx3Mh0+77U8ayR3Q
8pmpNPbbXYlXWsiWV5I0JvI++FnBKSNZaOCFDeSflM4UPTgHTRgWOF8A5d5KVktXdC5hrbPh831c
Dsy1O+nfuCAc6rtpdhOEzqNVbg84rUoor4/eosTDd212F07UxXJz1QcC/WKlIiuL/D5NFgF0dIfy
cbyHzIvLmBf7rwpJVkmwP9h9lG3kJByoQMXl9k9/L1M0mbUnd2T5TLDoiDVqKSLZ2zmWNFJSIGQN
PrJHQNnHZq8AYTAT6qtHxUNwra3+u+5dn6ecO3kKFNQGYoOf7fqPQCyxh5UTJbuX7R56xfm8HNSy
rNfLPz2q7Ss14KM6XP7Id9+3skOIRXIt6thTjqqT8XUbo+pVtZLk620enOYh4XIxqqL9hZA3bqHT
qlosFaAZNfGDoWCb23mHbhi9wk+JWGttZgmdTsmrbyDbkn7hU8Mo3lx5KdyxA7D8qipAfCxVxXhs
ifyDXlS38tGdzJuhPBkqumU0AYLbxtVYFIsvzqrZ80Uq7LHDPbmZvXEWSMAln85DvwZuXaBh2GEh
gnwKmkj6/y+iwlCJ+vQT9JF/6D8fqyCPC2fndzL4mMMFVc077AIA8I9KaUoFl2Ec21E19ajU9M1y
DGGyVQXkYe9I15+os0MnoNVIq6hn19m52CTvenwRu31j502j1RdFN2YYoNU03NmXv31oMkvCBxjH
lbUbMU0PnTt/6/3dq98prMxYMIsph05J4VrH0B5dGgjPVCuZ0uKrbw6iI94R8Crshfx7DcylVWW8
HC5oN9HJViSKi20nG4DnSN5bOCTgfIAXqBER2hB31bw9acQ4iNkWkIpIBurXersL0BK5iC7DFp3X
zqR4LLQZMnVcPvxoVuTEIJRl6P+jv0b4xUhewoGJ3m8aR1c9D9EAYfAqbZpV4YI6hPN75bdtevsJ
xrrfeKGSSOB5FeK7C76KwFlPiPhn3EJze1VHVRlt+b3wRsyQ2IioKPUXeZjAXIrRf+nmJnzo+C+Z
4/aT4+LNbKUuHvv/RNsDGsWJgyhYoqIbZZLWAB3/AqAYzHKDlNwc5p9LRwFHZsseSn8Zb+0374rk
xUXY1mcAe8eSY6gIJIVlVoO17KFWr+k2+ypOJafNXCwices/pDduY4DImHqf5yWx8d2ycvp5YJcz
WuqgSH84kewcr0bgt3aU+hQH81jJ10bNWCJsL4J782bVNtPMjkJRpaON+H6IY/T1zKfnAta1b1j5
wpfX/Dm81+i1wUVBOF0DtLD9I5XY8iDbEhwacZ2fsjTZreJ6rsX2wfNpPo7Oe4+75bISUHH1GKqz
fLBymEyYHSn2WMfcfnKPNtZldN3drvFU9EGoEZU5Nc7RFn5PBceM+hDTVIw48v01a9KH5QTKofNB
Vgk/JhLG/lYXapei+Ol1XF6OWAJKkRRt78tF16iks2a4j6HIQoXJ0iXZO23nC+B3GKJMwb3AKpRr
S4Akr/uQ+HvqD7ujHEbuHj+GevujJ0VsqQIvfCzprORyfoxHDdt3WTFd8Qup3h3bqlcAISPQiPda
WzgUeX2/Yd1w0+Xpf+W4rON9s+dUTrM1L10iMWPd4t0IQ3Co2M3v4PrNWdQYcth6eH5HQvgNPFRw
RWpTfD34b94JAnTKSmKBsnTVY5UP8ZH8ZuqHm50gAXSFUv3K/HGNRgIjlRJ5YXe4NPgXuw3VA1CB
xbTRsqt+ffa7dHS+6s9ClGCfFfxJMWp1WPOz3b4k0MAjRhTO3IXmG4EweKxMtCjIu8J7bREfE1Y/
84JewYqoI6c+aB2MfNrWgHvo2gmD+HLQIzYrBZTQmAEuEWYPstUvMDOAXULJC23P5b8UHg1N/sLE
4qN1ACU4SDCia/FVy8kiDGakNl7drKYSu7DoZafumVOMYzQDZa/+/mpPaXdfwMdqi01d/idK3DET
3N/kVmtE+XR3uDaTt4kU1zEnNHLvxOjaJ0YUFtipXVDxo//T1k1FjTycG8JFYcjeympEj8XBrM3W
j2SguOIA78pEFtuAduESy/qxClhFy09G56LxWdgYimdxnge8uuM/hgY6onPTMfYuDY7BPun1Eyee
ejqeHhWIM22lQQUKoVn5I2b8vv+Stk//YoDo31onIEBrQdB0+wVxpGosrqzma4G4Am7IaoP0FW1S
LuBKCy5BJt0P1PY8cbNGRJB9KQgXY7cBgua+xsteiDJIxU30F1QzaU6h9hkejjHbZ5SnCdRqbyvc
CL2ZXfV0wImOP4qBtBTIJjnk6HwR6Jz6680uKpVCHgEuBjmUWE+8JzudZAOu82uNNUTenP1Y9QgY
9Cv3bYjFNFR83TNG3ItmWazUhIn41CgkDQpEV5wF4lFh8NV8THuG4L3s9AvVCtoPaaT5l+YnURRU
OASmqUhksekrNPR52vPq4hGnEKQB34e1G3jqZps0a0mUEXpJnSeFwoRoyR7YAJEMxqOYAVK9DxdX
XqjBrrZHJlWUg00PNy2RP/HRI+7pXqgs8VApb8j11s1iT0JmvNx+WobViSo4odfkQKWPYYkwIqJl
Sdy7lYnfG+6qj/etjqjKDrskMGY2rN9xMLgv7NxSxu3uTWdkbpA1dPjoMzJQ8Qlka5csq8UCaxvq
zoTVcDDMG22kl7E3Kjvs7HfyH+WaTa1QZTkTNCRqU2J1Wnfv7fOcwiOupEMnuOeU0M7sYmlswyz5
1z38OKeZDSlKybxQUYl+A5LtgEUEVQ/Wd8zqa+lfXdHcpb63I6NoJw4D+VLZkdicLM/TyQ0KgeF7
8etsViIATDMQeEu+eiZzKWPh9rzBGNI8K2D+jMgbQ4pZsIxENdwJ6vDoRs2eUQ0Jd37X08+tY9h4
Hfc0k2pyKc6qW+ipC6h2R7b6KWH5JIdbJrnOV+cfGCyTmKRWbJMprwAXzDFB6rR2BL0lHRMyb+Mi
p+prchKy1RIAR4nND/jOICCds7v1c5ux5abGpMwS36qQKXmdwZxp85GHfcvzTvCVu4WxaRjKjLLp
n939ISV3Rgci3yqmu15eDOzWtw2HhvkoRzcQhuy7VYLPcA3NEZxEUNyX9lRFP6G8vwUv/vZvv8uW
QdZ7+Iov+zUdNgM1pI9qMceA7zZCO3gj6moZeEF+dYf6WBs72mZwi92SGWAv4wzWqVgWqFLwTFJv
i5b9Y5SLKX86pGpj5yMPGZ99TyP+J0w3uTVCFOnBTgIBuug+QbZtfzKdeZ4rZ+NL3/ZFcS5yWP90
ZZJIbbeZsLqGcLVZx68NlWMFnG1as6+rb5NDalPkLYjnCtOGBaA42dFXyLRgOjqsqRG+QYjtGbLc
kF9hxOkVQNxraOS6YM83T8w+8fOXhJ/gk1sTpno16hxXB8ujbShjsE4xgeRXD50HLfUc4LEqi/Zm
TzRjlCnG/6R3qMY3k2HEdLKw5WBbA1E8ojrje2NvVFur9siqh0o/+CW3ZI4peFodV/FQwIpSQ2cZ
f6ZksvnUOjdNV7vKVvPd1RbBLHqQLBmIeht33m9F9/xif4mvSrG3iKKU24iI9NPWyBNKquGPavdu
hU/YBt1wbPYqCVdKlIQFcl9aYuzC0JqS7AvfTqV4gD5bwVMaZ5CafsKo0DdyAO9ZJFxtH593VGe0
YRqN7aKFFUi17OGpYZadKZEpCBpb9GmiihigMwW8iSodsKuHX3IKdeZ6c9SrdDUUXmiRDoX+vTK3
pIP1Xmb/NLKfRslfPtF7TZLKhDX24XqxU9oVsLKuP6enNgIVyzVJBFexsSMrjJN9+G9JfM4kL1QX
+OvbdaOWuYrFaB2fqRfk8fjKoQ717bvglTy3BV8DPRhUqgsOIMgzd2m57uqoCP7u+4OV4kgQ8M/Z
jxgsRw1yn621bui/KYrqPiTxKS9TLMSYv96xJHp/rQsX3PxxYsTPrZj7UZfkMjomMfsY1/H7gT+v
xGPa2+96MCFuypp47iZqgmu23m9611VbTaTdqdwRKuB+Flrj8mmu824QRQbpknwr3y5SimjIdimw
MYMfNoFFjugY2R3/qP8Jgh/37dGvfMG9KsCyxK2SJx6aJCxcjfigPt+sxY0O+35B6WOkiJwh7Wv9
O/DSyT44MpZLHlHsIlk5yJGPyHs5vQ4tdtGAjpx74ojryhuERU1EJQnaS9Ik3rvYF9JPEGQhUnio
Y0WeU8sXQeDiJ0ICXt7WS0MKm3zO03aSMr6ssM67k+yBVEb7Cbz97T+0QLfx5ZdVpsCmGIIM9vz1
1uT3YVi+VlBqSXVLQrHTgKFk5xlr1Ibw81c1Afkv2dRjn3Jb7vVGt2AdmT5Lszbt8NRp56UNHaA2
+UxmRsysV48uGz3ez+ZmqomIabkgpimaDn49v3EVHx3KwjA+1PhMQ6j6fEBWchv5COcB9PhmP9tl
qJuILR/QWhjbNeiO1k9knL8kzybhTPxUk9e/klGXEY/rihWObAavh3yEVm4ZeFaFjZXZ7teuLosC
l4xnloxdDE+mkRBLgD9CagFT8ArQ/yE0sgP9oc+1Juo6+SHl0qqDaIa0LMrruCR+837WmWbYkRaD
0QnLnR4E9Y09rKJjTSpiGHRiY1lr7ddAUTMwQBDDW9dCCaoG2MxaVVo3YmjYCFXnBaP1maNjMcUt
gi2DVRm+ZGeJldX22T+N/DCpd72wW5d9owc6S+UUJmd+JX+tWQCsAIE4xwd2W/y8zJZP+eOQ/JSD
PYIOoNi03/d4Be3Hm3hpDYogz06GP72a9GEmKSMQs2IfLwwwdEQDlNCFxIvkn0Sb1uk2Pdsk/fdT
LTc9bdZrMuGDxMTjCaS6n7vhuYjdlR71uFydM8e0N4F1Gfj3sskzQwznF7ChfwmSrEjyxJTZpKnb
DWv/TY0CF9a65DdM6N4pBa9rgnWJKF0d/wnjYFGK3qE5nyufJs0qazHxQ3gBiRbg2cEJoneh1bUl
MdAci6GVL7R888ts9P83b3eqYt2WtcPenumS3EU6aztYhn0U3dui6qeVcTceGPrymyGcF2PGRHuf
Qi4yYS2rDR8AxJy3Yv/x1j3M3X4lZBXmxnqcLrVa8WtrNtQRHdIbryBtkRkf5o8ZYL6NNqwGjgfn
basnTdRePBvnF+bTTW6zFXQQ+fMeq7pahVeuFquIR7NZytkunUXJmPGwAZiLcxoKg7Tc0HNQYKXl
XtsoCGRZ6OLWBcFA+dvbbBAy7qny2cq++1bEzKmNHrq44BWzBg3yupbXPSq+YH3V6j4CcEBLE+BS
EwYXfw5M0OH/iT0JlCkBctq4FwbfBvKYxU6UDnu55BvU99M5t0F2xrLnz9oz5NFUk+E0kKQ6OzNU
h1cLJaOLDxJnOeXNdHnX1n1QPhFt08Z5P+T+9JzFyZWmMdmyp9KEYHaWi5O8vIazsWD/jLGasTaM
QNyJZK0KT9bwlArhF3XkZHTdoGtm6GuyMs2UfC8/E10hyMEF9PuUjNT5Omp6f0YxbDbMgpsRte66
zsSBo/OcJagoXQCs3pnA7ms3RvaiXABE2LziSROiNMmF9S/Ag9B/WR2qg0L7qZ9iZ6aJC+7buer4
ezCRcoKyozqfjDzCQBc1mf/iIGWb+U9jvtuxK3DZhafs75CMlty4L2f7RObdiKKJ2/BBenpi9wGi
cmDFEOwyl4pvlx/kOivHi0T2f/4fUjbq2qbZ4m+xm7dV1G5Wzu7RTfCeooR1U0ZzXOmB8pdB5zjP
wpOc1Feeqkk/fr3bqh7nq5zRQ0UbKcPw31xPXNNlIjfV/GKnceHV5ygRYKA9EFS/V44UEuy5asDd
uWFxUyTN1h6CjyNZWT9bSEY6vKsXHxyqcrkwnY5m25ciYrm2NZYODj5ql/vkfSl5PZZCA1v3cgsm
owhYCk0tHx73DkqyIKVc44++xZtPzYLNK9ZsVP81tWU4hgwTwzRL1nvTs/ki78gPNIrNmtPdGq96
MmI3cVlD7xacEgCYRIuRsCRFMsfDHI2rZSKYEoUMWN35WsT1985zboJxsrlacYNUaa6bozWaGBK9
xb9LAOhNS2cCn3fi7tP6YPRMV7d5RynqaIoY2n3r+9FOefZGBz+1O7gRV7m0iG+hX2y1VylIVYHQ
OMc/pFUnTQHcuEqdcoxo+DQFUiqi9/AhOryAHfHQGeqYHAq+teDQBnUT/k7+SQYMaf7owvTo1Jz2
BrqE7dKYq2iF2NygqFGPGUjb1twtrM/SN8XkGU1tempt2qN03zyyuK2sugeEoY9KjF/eKptEYTer
wuN5fB75Icbs7k36dvBYBnEubNFE3lunYliBAVgzUY2wPeBi7uVE9b5BZzWvPRbB2YmFpGXISlqk
K3WsNQmr6DYtc+gwyMLfBV00H3Ov2w0l6P2qIemw0QCVsTF6RFKSEUGmEYgCtJwaRCk27Wytmu08
poH9RP0/5vvhED6A3ggRxH5G7uwSeIeZe1xd1XPuk20jigz6n1e5PKBtgvan6z+jHlv0pR4yjCov
9sa98zW3vv9iIGWnuo0uszdaMoe9mdm+qdmBBifxF+F9IAuTrqaM3BoYeHxyPwP/GRNoD+Td/Xvw
SNcomAZ5x5jW3K+SqMWSXMLO8ZD7OcAjlk887vfOGxf9Ynkp/rcdHfEz6ph7NMjp1ObQzpkXeIMW
jVqPh8im55MNQ+0yW5o1qhidInSarW53SU+bGdq1kjxb8j8iy9AhXg8P/dNa2XSVLDLXNJTDmoc5
c32h9enGsWby2xKCIiS6qLhjFrNb+0vNm0j/co4AcCV/OA448vee53XssXTXAzUMVEd82Yyv1lcm
N/SWYwJYyKgaVPvdczJnMQbzylL4XvkGQOew61dikSMlR5HaV2q51EpGQabkEwvW52L6BsEgDoon
UyK3VNukwED064NdKB35QAbMK8eHeZeCfc/Z5jKtZyO9VAkrjO9Vqg44bDU2EfontmPT0gvRH465
UyEWGUDJOxe/Lpc+mh8bIODea3krLoohqQ34CLzL3dt9WRW8efAWUibrspcFUoVnbmML0sPwWQMB
/yAKj4+erNlcWwnrNDvJBNhZtJWpFuskOtKXkFfyvIdEwqjR57wZI/ApdpFFBhmu7aMCHT74LVI8
amWCM714PCJWgnGfjd7yvG5CHyAry1FwXibCOR/tEw881cOMS7iHbTfrgJqc9AXdkxCMdrFjK3g/
PAQhBIRsLbk/FPqkR/KCIzoQFbaqQZhW5A/BiSjBmXPpOuyouU0KKwDoG1zGIDdoANKZ0A0/G6Ai
MMN5g7XEAivWDxSMukWbBaPQPMblskm1/Q4IzKbCVUx7+3ctfLI/pDNBWm+yfDj2L8jm6AbJxuw5
4EQTz4LJhxOnDOSSvtE31dQjheAp7iaYirsspbxJ8KPwpZIvPcnHy90q3ntRz9PR4zsmMpkc63MD
VI8yWeYA9Dgo/2y2kvTybQQaBidZm4Nw4jJtJH9foKsbLbdi9/g6VAHI+oA5E0XCc6aU1rqVEimk
Nd6n4GdCOApDz2QNSYkst8uEiusTUAuycc6eL40V1+23G/mGpIhqS+rHtw96pssPdu0K6TA4FbWY
h5BjOk+2Er0IQR7NVFuZL0ZNp0WKU9luzoByr/DXZt/V7ca6sMEcH5CYsckEMpmGWWiC9bkCmvcG
9RCD7rvbNKy++CUHSoybnHYsi/07116lTvRYgi7mAE4flnBMaREMHC9EIwok48mADH0bjABs1HLk
vP2SsLKz48dCCrJ7vEv+kS2ksJxJRGkXfdSOtPfEp1MUbEbLcZIgAKNsmn7r3M3SOCpWw3oGlCrv
V8pJhqFV9q6WPruNfw7Nyg+RVo3gMuKL/d++yOXpSKOFLbwQJ5JLZ0fbYim5GEK955L2YSdAMo5h
IGUAuAAWOavd9hwQpl7ucht2QOOkHaJN0BiGvvuoAmqcl/RU0ES59kPm2MgrO/QAgiKMdh+rkkDn
MogZm+MEzRvYBuR8vfu2LvQHBNdGnqHU31ay326A+tc+JvTQOq/xJJ8fkmGXyUgkKsoYiY6jSNRp
nrxlRIeU20+jUunjxS+AzGlTfO2pUR3BHXRbreaWR9PWQXEYcq20ohJwI090rFMPqlxktn0mdnt/
6v5gefq1GDqm0AL82AzjAEv9s/W9tr78waAB7/zQ6o0iMrjI8PAUN335sXx9bzaCQ5meEXhsLtce
1rs2urtqbW9SO3fXgSuhB9cY/GUj3L7EyfONJuBx4dOUydBGW2mXmscE2FMg2DO+k0pLdsEAwgb1
TTAI6ZVsykFIEMncTJS70OidPRw7KkfR2VYlsIT7WvCuegUQwTywV0i9ol5Qa5WmLMvcI/pj1NGM
zy37PUylWwFTx2qBZvoBjuYslX8bwzR6R4dYCrRfIbhoDxejbaEx38KH8fUbYWX8NfzZYAM5Aq5V
HDPw2KrmS1FI1ESSavUUJKLVVBVF+S3/cP3eAciXQ4LQQc3CVIBm7e9bwnS1GrGx3rrFOvLhyt04
ZXuHZAEX1WaJbfjDAc9IXLcIvNnAZbd8PzSjVTeH0VbEGW+AlEuoxYZIKCwKNQSsSAjdIpen9Lbd
K0IBLtJLhrSrh9lYduCZL8lQjpuROF+wJ+yx4t23L9x9BccnsWX+3X1ASc6P2VeuE+ryh7vRjBId
DLsWIj9zqXLZitQjGND/6rDV4eMZVVQVbcGXQjyRR0Qys11gFv930Km3rJLY3jVKBKZiWl9WUNo0
KkZG68I0JhRDX2XQHcnfYBcTQgfY0d4vcWFnf+4u9pgr0PaGMhXnnM+KVloVQhDxQxR9quH7UI2S
LAWH+vWMGx6TolhR1xPKLAzJ4/KJ2c9/QbUjOpOCEk9ZFtLMX2vyt2F9WS6dGuqtrQ5D5bAoS8k3
B3McvoyTimBfbfwCv0anV3AHda+tz5IcdneU0CE9r2p+CSbBWsbjUk4eSx+zscSy6vjg6Tca5b/c
InyG3vV5/yMxUIMeDEX6gEaWbFc9i6yEn6UzMbbfwdXwsXuXwPVLlHmZHB4o0+q+gJx3b5k8bRxJ
vDtnSVb782UJkmrozvN5K+laNo1KiGA5RO91WsidOPiAFzO2dSVAmGaC/hp5qRIbgMjM1MxSK1fK
33POK8eJOOyIQPUelegyHcIKflIsn8TtPJt1Ugf6H0zNz+qxOq581Qiy1+ITHrxK1sES3L/xj6GX
vCp747pJEkVa/GnCUIo+UEKd54kJzT1S6VHTouZYOqeFogPwr0kblVrBFOfruCr1W1DOdLm6cmJZ
QOo40JAnq7haW5BlAvEP5Ji3PudInK6flTpyuolSlwciB+AzQEx9neFL2JNYqVff07MT9N2EmhFh
nmHU30AvgHLSGH13kJEK4UMRb79vLnbkgHnHSt4szY+oyindPBxzszwgy9sbSGpt6/3Pj7kXFz0u
JI7vjTl5XxvYSWKnBp6M2Y4N/oMVD70CXcCZPPc8/OYLyBXmhL8atPHx9M1+HbT1xdo8/2B6DfVu
LZodtPtCK1WZJIzEe4R2bIqZAYrTElYxybrpza5Rdr4mjVzYTVftZ7sWJln+Yds5TyfFi7HdDc4w
cEnqaTVOsSNQRtSprtrOfC+TA8xtelo9cgeGMSBsCLXnKRur341qgAaOU9EjEgaPoD6cvD6AP6uv
WPBtSnSFLEDoKAuYjlAf/yPEQh4SKVmHGyxJCt/HXi68rpzoahjzUB6tkYkwEDSL/Rh3OGdfY9Yy
UJ2iB0N7huQnit55gwR4qBJAvKLYy90u+OI2qB5DbjBAr286agNu5pKBc55JsBI1UjCvgTxOlsAL
ku7cGgsD5tf+Xyb2QXmXwMkz+OGJbkKb1oXovs//CALPNPIheIlMS7IOLsADof0La0Qz60FL8Qz2
AeSI6mPoUb+D/RGw7n+dkWIIoQc23WoUR+yfVI5WlraQJbHWAdcjGEctnSMSyGj2SRItluptHrlt
kjBxHpbNWitIBHis4PAOgLvK6FGfLVH8DBVUMei/JleSAnRoUU2rfQBV28Tgfy9AlyTrGnge6ErS
t/RWQ/ml9hwIMKyaoEIdnIMNx1l4j7C86DI/fRwdqwbBbv7D+u9Z4qlTXxAVmRA5MOSFf6v7piLL
7pp1wMskhDpVplNHdITqZtoP41lf+8vfKjIO0gXxxm9kfyc+ofOBI02GGBWO9LkY5KETodGYoz9n
mnbdbjHZHZEHFRiJHfZ3kSPlwIUtXJp6ks3YLD+7ra9yxLwLnPk77dZpN6jx5BpXywsDqmqV29dL
qx1k0kWb/wJA47WK3FQSdfETcoSWPvagkV3xP1Q02jmr5SmgWrod4EzG29DuAdO6gKvfgDBJoNkT
PTaLGTmn4KxhVrbxn8mr/psX1nSbu5lWLcys70pUyNav9WeS79LpScBaOMp8kzr0MFkBBGxexQ5Z
Qh6U60OQuiYZvTBNwoyPSQfRTXcsvD9suxGXCOtJAHUO3aBx7HnJxhH57hXNCTuC5qgJYT9xxBFP
7hZK7lo0Jl3+LxhONVgJjQG/NvOJebK80URlP5oIdub5Z3Grse+6AcJxLqXcIZhXcQKjgAZOv3n0
cY7PrOKDkY7a1v8Tg57PCqgTGfda+tx23QEDzPmkypikg9lhjEfKvV6FErSgZv5klrjz2FvPziR4
oBj6ygSqC73mfGJGpoxmMqKlPo2RqTXms3SV3WVknG6lS4+Shhffhn32U3vy3CKyp8+wYQ8rsOSg
Ve1gVbMQWQQ1yP7csJF/qQhs2oWji+CwahPupTdIO2QUkbfUY9ysj9AbHYc1vrNXJqmvBHdgJSFs
6XqoQJ+MTy/rZMOjjSgCspmJRSD6GVULKmBqQhhVDZeNGBMHukAq56VWaCioWFCvbUseoMPFUegs
9J+XbRTdH0gwovvONjt33gcf+NtD0/DFc+1ALxjjx4vXCMUgY/2wVdAReMqNjKSYsZ3/KNM6DGI/
mbcggFBPXHMA/ADps2df9M5f1YGgJBMsmef/fl+zBR6Y5TnogRJ41Zjn4/y80QYCOACNCjYGF5F/
yUtbVFTUzpcVOS396ytOyWa+3BnrRzfW1oPQDW1sjFwwIBb7ds1liF0S595ABcto/1MksUiNN1NV
sjGW/jq/2PJbX/ab+oD0Dh1YFGegm8cIrVw9BiPi6+5s0959v315+ARA2tic8KZ4VoEYpVA4q0Po
Y8CujgI+wmcHblELL1ij59xg3peTYe3cpzEsdkjWuEJBDQdjL2apEQs+NYe002esp987Vpg4VWSm
5d34Mk6kQAIWwhWrAC19B7To/PkrFzPohSowJmtzdiEN7T300myumAcSK5Jf1izc/mh/VMeBZocp
lVwATNanb1fWBZnsSKz+ycId7nHFN6v8hTU49umD+omm7njcKnVqMsAri4hHVFL8B1MG+Zd+rxNK
/wqlZaszRbB0tknvx1imk3s93NIFie2eucYNS3hDads6bO7KeWXezXDrJDB4wFV9lWnd3kYmsYFT
Kxaaqc6GBX1Lpeotv/+5Z17TRXqJjwQsQu+a8gewD/jVIOGJpKeXPGeHDy7R3PnJs3wCqD/MoHdm
MxjjKNtcQ93zTRrictaIFXw+soYR86iT9PnMP5ms8c6Vrii5s4W+JeI46pSWrQTu5N4CjmM5zxDb
8QrASOC84c2Xp7pzyM0uzYC075WuCJV1UBmAQy9lIOCz+38C3CrAbHJFiE7oi0nJpzz9F7lZC/l0
jmT5ZwN1AnTDeZZEtBUhNNQRnzbAhId3f5ajp9VFeJOvTjbgMbsFUdwwDjUByAqaLXOjj1Md7iMZ
jqXj/pMdtjwOjra9sLxREtnuj1eLcwLEQ4GnsAS2w1QdUoQc32mBF0W+eGt8lDWentM0hDlm7BvE
OTDZpDHfes0P32WCEs1xEZ+JKLdzDLswkEy72lMUHpPa1nETM137imMsIHY0Iq++mQ9mY39y6veS
oEQfs62xl7TXCxtV8pE0ZzGAWz+DikvMvyGXOh/xGWXZLW/0UC+amqaRjE9mBrA2zKww07hCfkem
/dwxM2x0fUDYvky0pMN3XB0Nr+KyGf5UPKeoQHUDOMds9vKlRrUbIw2IIqCdnjQZSCgLgziLqhkk
9LN6Rc7U5A23dDH5Wv+aL+YhRk7z8vv6U0ghomiyLJpR553qjBxQj0I2ezpPYw1DfHdgWYVYIjrs
RRPvRpYabbVBW3xXDUCdUGZDrH3QStHcqm/dfuZ7OCHuwwxSS4GGr4J+2rBYVImCNsg1NQmlgBsE
EIIUfSLj5VAZrhd0n3+iLzGzHyOy0zRRcwBZYJp7jNeBgIyZDToS1oYZqzapPwWLA/yA0pl6gZsE
cbhWm+oEazJY7p2aWeo2WH8CY6jZPbqkwtUTzknTZEuEeS3INZwZ9TNezxZwjSkDIgfp7HSJtkLQ
Hje0zdfTS4La/mcy9QahlNNe74r+lQuThDi9/LHJzfyGMzeB3d8MVc2yqfO7oR27Pgd9Gjy75EEC
tTm+OnMkuz1oYbcdQr5P0RlgSpWsxWAOhwbiFUEh7yvkl8TP+Rr/phEPEegklDFfZuD3Pocn0cIE
Ag4fR+S2QHgjDxUcUac25XdOhobrq2Ugi/hu05SbmzC5lI76lt6e6mUO/UZD96XXuGdOZDjr6XAG
12DYfTWrU10JPaR14WJ5KderamxMgDN/1qmYm18on6dtNgbp3JaktdAH9qSpeZxXlVPt9rgKukDD
afBJekSu/ttxh+l8ndcRpzXV9vUaAwVfje63XGyrplnu5NehhRlMpXj4QKAWZ46tyfAnhWQCO9Lj
YB8XpNzwhmPugUhiyG9mDMk12T2omE7YJ6Os4aJLiGCAf/ExMTY6GKWfWzfdAbGO/4aXLUg5sbfw
CaqOpjNho0wpLN69JloLsEew/l96i0MVGkdMzk9Cfk1uR7RSAIW66m1TUWPyfdfN8uWxR8REXz4x
kOLp3qX0nwRZSXdtOuRsBs4zKmwlIsQlrSKBtKrDpyxPVjNBjeK1uxkgBMkKKNCHX4PUwePXyXLN
It1vsOqJfDI6Hwla5+KdmR6rzk8dBPP+X3e+rDxdoBnQDm5QN+xg3ifOb4/zRA1QNzIWPZRhId7m
AJVqs0oAVHoQQChJk9Kyk6PBfEWNdpkYfk7eejxbWLUOZKwWOOzopdyyIdFsg233cD9cSLPJQFDL
OyWix+Qxz0SQflyMU2eFWu24+L5ZhpFWp50nr8zo36cIU07GVpogCZu0p938hBH0JvllFgqDacqM
mapD3LBvS8gdslEZzjC+fRn8pOVBCL9ZjPAppwBcaZQPHwINGWL5ahGrQukgt/r6ZGOq/pGGSxDZ
sHtbA+qsU3gdpNUlTSsusmCtXLN/tTtiJIFbB91xirE57ycJat1CiP7+a4pi7Cpp4a17vslTYpXJ
diyQzwnVrZHaW08nAnZCQf4OyU8ntX7K0YRnbuN1fP4GdbgX6/UFN5LRyM3Sq4UZypTcjqo96yQV
Ucal4xFBaPoz61w0/weL7PVccfXhXQG5GYqgu6PGEsdL3o4I1wTNsof41crdiyU9zo+d7SGZ62Nh
hDuR+cyyyjsGBm/HHMLqhpCMAh9xze6lRXphRqSPVPoN3ZoDNb0xCjeL+UjYH9CsvFeqGffAK8b+
Pvux61aXQtwFmdj3BDgNn2Yv3HBE+8tCSeKHk6hXDaXRowk5GClp3czKGmO2YmABuwUNUVaVp+St
UtdIJ83qXARRu8Od9PJ3WBf6ZV5ChHWEudhd1bhRvOuldU6FDT5kOW1G/B5/mH/IuIsCJd/9pQaY
TqHqPgd/uZEbG4elRVe9y5MpizJSDkAZtyDXjOM2sFIcEhmFD9VdbN29i1pm9peJtj8RIWHPKA99
WUuvv4j2OklscNXPOSlug7R40T7HbkbJDeCbnNH3JG/DfoEOTUoRgyFNns6ZZ3tU11CsxFBVJMY+
b4HVfpkknM6ARZLRZtm1wIUjGyMvRPheATa67CWTHwjzG3jM8VQsGrv72NdFgKMpWZ5grK+P3gSS
MrfK6l0c7C9SVltVr4pks5ox1fBb4sPkxKWgmmhaMBWscyBW6WSFsMz+WkrtWbH8fnZNNzg30vEW
+FJzkmoXBa/pwq2ClKWDqTVJ0wZxRd0D40SlcRkV/O2ErxZoYyETOqXZO5ftqMGs2Db5FfVzmUa+
UcZaQgqjHlsGUa8fNOXxWpaqrNYI1jSNgCiYkglGgCwTCM2IGBAaI6x7BhTtPeAzyO/GJkTvT5bB
CPWuL2X7Ve3+2tuS+YhCVk8yjgWhPmzbJ8dBtyZFBM7OzD4VBGHJVgD3LbbdijjkrP0mtdVleTKZ
fnssoiAmcboNXWSlw2MHsbwfecSHTGOgyw/Uga0h+1NPlpPiQLaWbTtwZ/0C3XLLG2r2cWdSkoFK
kUlEYBwR8KtD+LmodQ/+fuze0v/GRKycK5I4DnwJ5mBRZ19Pt8vIO/ww1+SeaON4q8TU25G9GS1R
3wtZJYtMcDcGzk1Yt9Lu/Oumo+uBTcimP7fhUL57J3epBA5Mbsfi8k1TnUu15dCJ6HPwSKWE9olI
ww0F7U0Vpndxt1thR8hcfb3MsP9bag8/Xr7yv5C1j9veJ4rRpZFlbdEnGFFn+Q20DRFgGu2VGGRc
7wVdIuS8icV3ZokvgsrpXryEUsGn0kjK/rqwZ10B6LduYOkKEDLJLeBwz6kerylB7BcvmIQCj1N1
HCJ/2lvOXe81MSc1iL/wSD3202VV6mwbu+a600j4H8EkJotHpkirOmz1ritBDHezpby4EfOwT7l8
4jSyV3QDXjZE+Js6lNODwvdvpyHKsjUNOYlR4OL+iYP5uiHPO72lOpRYTfWkLsCCjXgVuuwxWzyZ
meR8cjGh4Hf7cyc4SdUhR2mKmEYut7Kg/ov2A+Zfrgcv1C4UO/ABGoQfbdy+qtPSc2Hdsw51pO5W
jdUrd2MCpiDd2ziByDjUX767VoRrznnJx3Yj2YRF35SgD2v6idhBR8rYU/pTZyWhWFd+yb5MlIS0
pWYG5rlCtiDunYRi8xyMGvLHDVzFAOjx2usB4/ojCcKSZiNSCdytNlRFhNuuPCai4Eq3mzdZFcxg
Cn98G2IcYr30NiBqXZCCH4jiQ5/vmstGSN04WAtskkSv0F+mOkzIDiXPBJsKYaC/kKLJduNrdBYN
u/czbaqOQGVz3LGmW87wKBXGwtOK9p8vkLYViGlQg+FrDigEmrCnbVfbwFnxA3WP0wEi0mAekEKR
R2myX1pfBX1/tENs95vJvY+vho8Mmo+SsidP3pCMDFKLJ8qIMqGE2CC40ounzo8yrAdKPahpfpfH
bAuRlSqmKt6Velq5fTj4jJssSJ00lFWyJHcqyT2y+/nj0CFy11aTY+yGLl7HISACvkIwC93ehOYW
2FxtoQqB+CnI7TQ6W4iMA2fOuZ2Kk3LJd1o04rfC/qI84d6SxBT7Df1F/ph4TZ2vrb+yAX/+t4ZI
Pck1mrscOSE/oWI3Xzd7smG6/EsMPszBIDpcDzHpQtnv8vRPTMWbyeJbYaQkq8dqOMvKos2m8hKG
0ZA86OMUAzigjcQTpMmpGLQF+KRIbQF74QgiFQRNItsd6I6B82cTVzAiwnmk6zwozT3NZ29VDknU
EOyNgMHQ4ONMM0FJpq4qr8tK1Tj/ZeXE12UvXO0Vma23L6WnOCfICKpcjt0eVVErzvDlVNjXOPq8
Bnvg/i9e25tGPkvwfafs2u5l+kTctiBZPEfQUsS9QMF10m/FBj1tMz/mPIN/OHNRvQx8M/bBszJZ
HqVuTCQpK7MibE9R8prRoVK09f+/GgBWxdI8pcmty31xZt16DLfGkMhBo2B3BdryzYLWk5Ob9nYp
ZfuVQE9tg195C3eAtEeUKRHlNp81UsDMZi9e+TzO12zOTzpKSlirGHnoXiKbLVb6mr6p5riPNZeY
fvA96ojQCfH5ce8wRAzKH6a+0RlltbqTCTcS10b+/TUYvVV546c/mZIlFw85CwbpOlouojfKi9uW
0O4EQMd2aP2jaqnfQ4PJyT/d3c7MTP61ZA7jPE59M+t1vrFGW3sXZNF8WUSE0vTAFUlw+fuJ1P4Z
UwjldXqW3fa4bJnTlgRr8CccJF3fpxm4KdEhtghkYs3q125exyAhCONKuFzEDD4M3VFHuA/Gi7Il
kdR5Y5rhoulBOep6dvIGf8uWNbb+gSxwbENJmWZSTdPBW4Etdgjj9+9LLr9QRS5/9Oq/BISi/5jx
0oWHwQ91Xf2S0oapcAAgI48I/IrlWlGtksGYvOgH+X6EL/ueBeRxvH112UX2m46OX/Qg/N1eWini
Nobe4wSm/PbVxkHQnR89s0Qg/Z0yXZnZiPjpZC9V5VSwTDh6X77kYkxQAXYHKivXqw/CWhvvtNgv
ZDH9geCwVKxzR+DPVMaDSfRIdGeMWFWjTRYN7X85gT/q//a/qOpdwV+pnhWMhuTf2aFZh2GxNO2w
zjQkFeEdStr45z8yEyBeZh1WdrYFI8Pch32yjloBLSzfXraGVVucS/w9CFqo/CEv2+3JyRAxCTE5
Q7mF6Oqr0qFXr/MoT8l1EQJHvQsz8EOOURDP+cRZN92ChuJ2UF2nKGbKHdChw751A4CSDpaYtdvJ
bJapMFoziDdROKi5mOwn16xEhkB+LBM/PqMhktKY7V/oYDpbtPDV8KUaU+DpWuwtNSHRGwVXHraE
3ORo2EXtqb4l3AgAZGsMHx9/dDLMpVACcI0rue1qOMJYoPFvMvY618P+vfaEUNU03kQAUFHLRQqB
lB1lPO2M1cWBJeXIl98kLasSHhQGzJoEMDovHeUI4+yZYX4PkZyDmI9xfIbVhIex25tnVXtPf0Fc
Dm6oVDk+TQbme/LVEvaW5Q3biQhg+Pj9yTY2LO9QN/2CTC7lNLK4WwakJr4C985i3lOjFBavudGV
G4KM2WOSMZ6qvVHNfT8GV/FTUuSpMLZavPbPIWt4AYKn0wQ60UZB+tPdxzSXK2I3mQq/jYqO9JLa
D3Jam9wh7IJqR4gTGiib4btC5PamCz0KBjbv8p9ntrMkgsxMU5yvm4rUE7TFFwkVBogG4XvSRBW8
1X5iAs9Ydc1pBHfeO+8tlRvo5RB0m7AbOm1tZnfbmjU6mk3N/2R2IkIHw6VS7mSVgHjYpWOZuwpE
+CSsXI9VKub7ySWeq5L1mDkXaxey0AWE+rPRHB7+jduSZRux4AROM0eow7cCBXr5kwtRjUeXvF+w
mc2rd9rDE9Bg+qJe5lL2VPh5u4dcBJOmcP37fVnTCXXZMwawoq+7Jodt1bDOAing86hgLj9zqJoj
Fk7EL8Duv8c4A5a9/e5Lmt0yQj4jocueCwwaeFXFv/zjo1IOpJfpP2Iq/LvYCHaY1/jEa5qT63lP
eSpDtlp8GJuF769qj1qUbRXo1D8V6G5qRjZFpXxvYxRkW4egD4Lfh8XT0Er7ysikLNaF9kHojfUh
g4Yma5e8LnW8zo4CsbzHYJi2BzX1g9ZcrQIUgJIO/cBBbYFTS8KoIejABQEf/sqFNxATaZ4lFtUJ
qkfYHLEeSyQ+Ju8V8hX9E7NUN+qwFJ5PgqNI921ze+c0DFfjHkg3+ti4FOPKmveUjkm9pjSAzCEi
+rYeXF+rVvJ/LzlCv9920mCjz2VSf5N9Ej/Rv3LiVyvvhkdDGGY7zOd2drye2CR+ewMhzuS/ugcS
j5BkRRBlTBW0QWxerLDh0MjF6y5xvLxgfW7JHRWf+RsiIfmkiU7cPWeaqX2SljPeIylbrq56ogF/
V+BX3I/88Ymq+sqDgZn8uiuvB0gSZHJKFa6DIbXNah/f+0OGVBzd1Afj6riSV2PzQhRWOp4fyvhy
Du5KE8njAHyS7sa0TFGgp6XhrpW2UjbJF8NTKWLNNFQ5L9FEaDVu8xQS3SqrZQWiDrwmXClBrVql
SurD4unj0tHERtQICWbHSYYIEAMVYoLwOe0VYwJt6NzGO5UD0H9lrbWGLXti7pSy1P5WPvNgsQw/
bZ1uoSawBJnIAgKRagM3xrMx5ziUKAqns67hwVgGoUMEYRTQ/b4f0mWFvl4kTi/cRHPfw8Oxwouo
F8qwaj2WexZWVzd1bE6+T1RuhLPDtCBAqXgIaAUlmjFmZwTlILOuGIH8fK9UDDpUfB5TDzpg4K7h
yqyYk9qhRPNtFBXUoKZrv9YnNhBhU5D5p/JgCR31ZDIUhDvljEp/oFkkhFxRiAAhb2Kg2qcT1Yco
mIrTDo2rBUNBguMY6o3hSB616DOHRgsYLbaoXO+EhpHdUk+uI0ZhX4dR8opA25/RCF0JWdZw1pRJ
xI35IjVV31S5LQMWhHxyYdzbGYRADU5dYiZUPDcq20bASc4Db9Y6Pmcu1gTug/MNW+7dNowIcnbd
RvYSHRDSTlQnqpD063YqS0hIHmYaLMbprZoCSr18yRcB7yMi5e51deHiN2lpIxlWTB+1qheyv0qq
y0bLzaWz023wNfKnYlm09JDmCAgq1vkeg8PO1nnYBNZNfX0FqVo7ZIHIgR1tcVWXv+FThdRIbf0b
jBF1Zu/IvhixeBxolVX7IToNiPfdo6j0a5ERvcPWDJv340dT1wCnYfiA+2V0ftAl41p8pUYG4NzT
5gXwvlF8vWgpSdRnueokGR9pZH6fwj+smUC5+dmytOsVE4lrPsnnQFJy3MO+zW4QzIFo6VHRGGar
9pWYj0Gt8ZLsr7wORY27fepPb1LwZh5vbHvg5iL1l4TH70+ZA4w5/Xq+5gdyKh1iHr7eipT93xGC
xx20H6s81xm0Sg/NXkG3iZDdkdhFV0emCvuAkPAmIeIwf8/6AEOsst7BMGGvgZ0gzL7Dxg92p8ok
+a8ayE8vdd5UEEKFXL4dCRaGzTaYSW52/Thf3Ot3i3yNb2k/CljrosXlqESaFTqRB+mYyplvcohQ
BYoVKf1xe3FeUPLXEIDGt+vL2QK6g2k0NSF5dNNvrGPtqqQ87MKLNH+Kk5cwijDlgQRfFXDQaeyk
vIAh73hd/mclC1xpTYZtR/Yh737VzLv2UT/oqrG2kD+DpEuQhw+J4V9ybp74FC6SDTx6jYakam4H
zo1LY3EzC2tp+miEp/P6ANQYjxpVZpGqyOmSaxYEHwMMu7NijKRGztciLq/vgWTHw5kM26qgfRuk
rt7mWHVNvck7NTj8SXAg9n7wbYYxfznA0NeByNRvxmu+VZLAbInLsaUai7oSJDKtFafeyFgzpynF
GwPLRj1zxOvz08one1LcmFS7JxF2G5zNR0TUfmDdxkBEYAeRsiz3Sz3zzTHb+eHJ92JHICY0jw8m
+kWo4YC5M2YC9oepptQOoB72uvKHf2tB3G06T38X/2vvPCRu0wzvjfEzcIHEhI160qwqgy7+yKCI
/mJijm7HHCYvwsf++zFjt1PcK/M5vp2GL9PB4winzshafgl+mGqkDz6TX+Vrjz5BvhqdodxFyZ+s
kHfJ8utr/RJT3M023LpVW5+uWDf5VI/JDSE62oLh8S0c1htM3S5DoGBq7OPaqroWFof1QBVkebMR
SXrsFK74VEAM+wmzSXUpLB90gRKjNtYjYl9tSCFn85BzHzlccy43D5uEqHgPHwZ+vxiU1wc13FI3
07M5WIdecmbKTHEkm/w/Qo3OO7lwbJanpa+gSFAKAI4XXZEI7udXucX0N09hHcY5WTpVCmXWlwGR
AlDIBVtnN/oAC27+c7g0IXpq5ehIGsnywlmMU2LsRhojn6tfrsGJoAa5N+hASP+G/nMRAjmjrrZy
M4YRK6nZGqcdv2Nft2yYhIzeh4bueG40GvVR6NpnrOOCTk+HioDB0DwH6n4VMXR/ROXgguU4kl7P
zZiYoEHPKeWBLsKRp+RyNPRMml48/ROdgN5R27GX/Tz0AxvI+2soRYMpLzixsY6f+b+PvlpI8SGk
t0A6vfKnViKts+bkT4ABVjk9UumJULvgCVM/dJ1i/nsv0lbhe+PLnjnGObVwQlx/OfkIUh05NwxV
WmjIv3/Hc6Lve0m3jXI6woxxH0XuSk4gbcvPpAQhu7Rz2uQO3esdPNySrxToqJDY5XYgGIE83Jux
gU/J9cTKOAaDzi93OWIhPBcgeTKuRcNWTR/nG4amkQToaxiJLauWN7fNoomvnfNoGKvCD/beBQ58
pHbx9h0xmn48Kp2iNs2B2ryGoD8MC9t7hLfJ5QDIUT9okcJo2X6T0fBKdBTcc35CoWvGiiMw2JvE
o2T3oofAsGyzWgOJbVXcFO/mDgwo1WZpvI1JGVOQ2C9QHxzcxwu5owr1dDmhd6BDlr52f8mnx+bP
PckowodCmS9YBNkLPThDRn0RGYBMK18A2KiVeUD+jugNdkav5iiWK6LYrhfpislZWHIm6F83DZXk
UY51zpWu8JkzJIEk2FxZ/mvWlGj8306NGDfd3KWdUoazv8rfVsaB+JpioHoVBxs3Sh4w05X26gjC
vH2K+sOpnwirPieavoAQtugqkq3H2muZLEVGfAkwilUcX1/uV0qF1nHOaKhaCtjAWDxmB0tSHq+3
snkU/WjZkMDMbY29gdyI1wbE1Lc/RaB3ClcSxTOlinj/Gihbp+Qr/8yoBerE+m7urIZe/8yvlw3j
0+PZUlc4mh6dwwgOko/580VKyHG31hnRuKpZrpI1GlQjzMcHfqA/Gn2V6iZeVIKufI9Q5PtOlJDV
vQQMHW4N8rr24ABiMO1EQVOy2V95wD2a6b4YcOj3ecM6GqAV75PiL8OG+f5durECe1gUi5ATb7+/
M4f5rXizIrGHvC5/5/3A6Y2CaALQZHzOnghj4yqP171ZbJJDVZv9+IYiP88b/dFbA1rJX04Z1u1x
NC/mdgBhgwFzCY9ZG4Iz05MQSjuQkJaimdvXrsSe2Bz0kCeG88YvwDumcWN8ag8Hk50z7ftDl93m
q3RPlBDbyrNEiCAjKLNzDgjMHJQUsxVSqdoHqiYd8B7eeyMAtQHEsmXYrKnY3zlquAjeEa9gtVXa
Gs2A5durrrWStFgVJfP6X1/Dd/fjLqaYami27mC45UTY5W/eV68cv6LupPAF+2C86oFrly7/PGp3
uEatDLgFBTho5Dc4Q0/aX8ZOBJtkMkON+JvHSSbWsy7HCkxf4L/KxmvEgJrrlgR66icTYFYWuUs5
pDHlMWG3s8t8ekc6qGDcYCGUROGL0Q1BGuytzBJ7WVKmOOBV8wO1Vy/xjwZO3O+DXTp2WMekLAjx
VpRcd69uVrzOJ3sq/vSXAIvRJYfK1tjNnukM24mc/g41Qa1P98xRGNoRu2KOWM1mmqssAaMdfPr7
MkuUEvhDNvWHySRWd0kWZX/g8v4EIpz177rm7BjFQ2YKnx53QyDGkL1d2Q6LAI1jVd7hTh+9e6ga
Z2/7ePdd28tQ8yE/rbLI6p39jn0qfg9TuPdHgeig5etyC3igDTLEBnDh6YQ/HqTek3Ma7UP5nZR6
RfZ359ThephOI/gvp2o5SeI0UxJmQE9xzQsJYcP0S5zmiN4WwGHkFkMIc1Tv2Ukc5sebRRjg1Mt5
ox4T4k6CMmD62AA8ZX7TZtbb3mYhfB/otMN3JTuLk3GwFtJUWcAs3XscUwxi9BOj/KeqwGURoFcY
xspC7dgPNTtOJzbasr2x6jgiKpXHrDwmd1ugEXA/eReHAsiiemHl1h3xWvMgYHoQ/oAs/wDpsCoz
sRhWsBcLu2GOPFZQr8B02kyxvoLgn+Hw8riC4Z+d587ncnPcghn2CMuU2qLaQG1mTznQr/WRF8YI
JAVbaiEeHM2Q8TS0rXTx76kNCTFHY8drLqNRafk1UMYSIQgxryrd1yyro1gWlKf9HFyMvs+mzjzv
WV5W5ewpjewHxGsKQkPQwJXx6mW5apDAkkO2AMrEZPs/F4JhJ1DgCUJEaudr1E/lnmkat58X98Ji
YgvxKOftv0BeR4sznFS6mwNOgKThftV/BiOK3oImmZjnyePtjnacFfW6m9QKzR+L5w/VIpf5+RT6
JoInQ/+8cy+gw/VM3+CSsKsz5I1DPrdMHolb4RkrtRp2KJ9sfhWtGwytvkhx0i3nekXloYgQbrtV
96c4wVUIIktBLhVDtYHeip0o9NZG6Akq1tzMwe6Zpo6ABPnY6VAN6iZmZZ2f5Dp5+3YQQUIHwfIr
NAo8x/7nDArFH1FBWZJ8Bo4VeHKSLvhaUiGr12eXdQUY6hoouabIqYJ/lr/+2ZDul14MNiM01uwL
e4Rh5L85anV0CwWkuwAm5CXadg+N2YqMw0kwYrSezPeb4pZWfn0/rYwKKrutvPWjDHaZJiCyqnDY
ESE5TOvjQyTJ6lFxElWt8WFYR//mvh8XI0GvPQSWAUQwg1SkHZaapRuryQyKPo5CQXL8GlHmvi2w
GmWV+pP4qdUbs9zXGvBN/m1e4STzSGCnxsozx5FqEYPCJ/zcWO2+cqpm2vX1Rd7WEpK5asxRXXmt
DdqYI2s4ir0jydaA/UnnHbQY3yi1C2SHs3rD79GahdUDH/0GbvLbM9z7WJsaq22b3/2PVU2m926r
e3ndwyOZQGwzKkX0u5mgQu5S2fxLHqbE1icqf48hKxtFdM8P0CTplJzcWkMhHbjamfaSEt0MDnqg
GwGJAE7WdRB7C5FI0/UhJ+dE/lxHccmPikZ/l4WKvWV8dE8DWVmDcpFqKQgGfwhU+My/4xbrV7Q2
KiHyXqE5VrHkevU8lGvkPxJub6/T73g2BAiL2HjgpBL6UimVyXoax0Wwoeh6XSLm2NcWvhrsKVw0
4unMSjvXmLrDyWmJeCMPiumGxlcmhG5iyfNCcIEr5MLFERT/04zun4CxRk9mupYFkgw68t8geLXa
D7c6HZz/xw5EGXba7jEh5EWqFwwgb3FE0hxYzjhFNYq7wCuEH2EvFSk9K2Og4KRNs9yeb18Ar3vR
w8Bku2S9L8hS5t8I2lPRciQblBy7ZYBTdIo9yWwH6lXOA2XC5VH1bhgCRQTY4fx4OBnTmoXQPrX4
F9IH0VYkUzlW1JoGPdqGHzPCUf+1OPetMYKGrq+GJT26q3WWXi5svyRwtMvKQOxkStOzEjp1ViUq
Rwt/AemSfPlRevSO/sZRVbR846Av4qADE/Tgcf+1P93VYGS4siUyxQdFVuI84ZhyIR6PQVN78xSS
D4Br95g/w6MJf8tOEEeDTZZEUhSRlvbCS29IDBnSPxZaumHW/uKnvg4pbqk0u/h9zX7MYhYel8Wg
rkHLO7q435ZWvlc7yas3mKdshUeXU+bALR1SirUpARIGQDpT1tof4I1wMp7nZmUA1zut7VYFQXlk
UOeGNRsUyA3G4AsCnYRXHxDWW6JoQa4zQVeJDrNWk4G5GqLzUVycBAvnWrbYyRbDPlVzVnpSGGeb
WM84k9WxSdSIwDBodk7HqXPAz3beWNxB9XqapaEV7LeEcZJ7PdJo97lTHIYThWoFoS5HjWtpmbBi
ot8jx3FUgC12rWqwc+jJXkJkr8hndX8VpbtC+LTfnmE+c+jrCelbDbEOaY0kEUQqQy8nP73jAHy6
h4A7MKe2ipxqf3BU9Z+1kfsCYx1pUTLLlGvoxegJcx4fmjiTGDxTsV8a9RFhcv1BLCBR+nmn+NYL
SuTEbNEUwbqvwng1V+y4Hya5SRm8mROWwa/sC0Er04HuSdoQgY5PTFjyBOx4Gab4S4X89bMnTaiy
JmruS12aozd3JYYoLsSdkdsyEZntV0ZDBAJ8NibjQLiHPtdVgHcugh6QLQ4KpQUav8yR/d9ZJITN
v5Qm9rZikLmixSgh+hJI9Ob1YyZUyPG+9a1WwHk6P3EJfQOv7+FWRvB0lj2fadyT10Iub14T0C/n
svJ6YMmhoWK9dczCJKS9Q71e9wgo4SGXlYXBTyy7wK4jlMlrhAjr8UU2VFXAoYyVEpAroDbZzBoa
ty6ADsGjJDaS7Mr873sxG8wHwH5Xdx8LpZinhgIF6cgnRF08PwEF1kNxtV3u0grNcxp4qRALRt3o
XLGuiyKweTpV7S+p9Z8BmIHFqG8vPi6B2oD0dVTBZpgeLjW34krktn+KXBBednNprwOSqyvgta+n
p36HbYUzW/vXGZXlhZCTcAnVMxWFfELogxV3JvE+OCFTZspdHTL2l9U6qyp4GlW/wHWs4IaL3CdU
4qPnJ8eCWHxzvIIo0RIAg4o9D5m72Uc1NQZlMhoHkTQGtwYVTO95jXC9kLbVP6VpD3NOQTXyhRbs
xwOQP2eRXrxv1VeL3lqh0oYaBWaU/RHSg1UbIjZdAWUA/nP2BiAsH1OVuxfCO58bDRQAR2oRze4g
slyrXW/udpXAxikttrGVQl2dgzcx1oVBPf0R7+Dn7NdDJo7UqpsKt2Ex1prqjzddrmdQWzSjOpQA
c7nXDNLF89FBIK3TSxEvtXqGkyAAccrPqEwWs4+vfwFkQNp/PA92+S9ojpqXzx/BQgQ1i3bqT5Qt
YlyEDIjOfIKBnksi++4AkdeqrtgxCXdhWyjEU+yqsjdhhFRdQMKclV6whP0jHgHJFxK0Oh6Ovnx2
hpneqpL0GUrzkrTBatOglJuyp6Wg5iWqZEvnPRpr7oFgLB4jftm2rNdwe+9TByHs8+gCuojT/rQt
XrFeWKyfQdsYfhnCYCb0IcG2zM3f9sWBqnYEKJ1VJJUVdO6aztfiTYoTbJKCiOXwAkMtFTiX5zGU
jbrPvZymTmSvPTZQRLY6Q/LsXM/9sT5gw5j0IsQ/ti5Z2t/rEZXeeQwGPjEdN+ygC4pwmQZmJ9yr
fyL3ljqZ4Uv+JvTmXmQsetKhJTBw5cQUFPJi4hFtWF1P8KpMwfPj8R5IIOKvLLGui0TIuivSDHkT
uiofZdtujmoAlXS1pY8GVWUAXRCfT87oJJ66X35VygcFEdII4eXRS3zzha4CxIFMRHN+hSt5W20e
CDnJ/zpeRrvEqH9uDSkBsrcjNi5xZDbBlGkcXGm38c25qkGcX3MCHPKPVIPWGm5t6UYe2Tt8ONhX
Kzy9kjLZGJAWqJ+L/NZ9zOuZichbt+8H2ZA/GPRzomZwawPHBo6uSlc9pxkv1sk/UJe4LzquaBU8
YvkD3aQNWUilh6LvIHOLXKq794VfLSe8ghUeKmOZpLJ8GXDO92QpB8DojLQftj1uRfPjCRYlhs7y
NOGakRU/QAOVyfr1keE/NOms8uZEg4Mg4GX2P/KmLN+fkbbUV6YZO/oy9BUaBy+mr2yr5zDjIryH
Dnxa2Ri0hz8py8kvfShRM/DjK0nYJnY3Mh4ZdGSl0giDbcD2MOUQLeTdo6Ks6QysamOa3XT5BVFi
E+Vp0ZEsVBYl+BM0qs15/Rmhd5fEb7UxocWfdKnR30LbQ3o4F+Dljr075VWOHztkLm4w0q8uqHyk
jamqoidjJgkGPKC7C6kVY9sjP/6M18RE6lmgaAdDAxjGAfZdoI/3Fw6Fziw39N1uywDQKCxec+Ri
VQNyDZRFLdb2pyMHWqfLzq3LkSejxVohw9t6iBmuqdXtAuvjmS3KdaRk15N8HLkGQWoMpinxv/o1
rsman2X4PnPYLlRUCWMFLpLhJTMvXAIABekP6+orYGlesVYL4M3pC+x0vko+kMEG8i38hUBx8cLz
R8FtRUI3V0Ms7vDrHuzUyeOP9wtisuCRjZgBjBSO2ZcU2eblWINpn9dLvKGxB/miw9qdhhecIXSy
13OeItX3LCUT+aPDUiYn5miYI/s71T/zUpkBAAfwhXJB5GCQoGnHxUVOiMstCm0f037fV5T9SlyO
f+fc0h6iLxFcbNphYDnRfBaCzW1Rr4f40HMuCkJeVguSvuTc2FvIVLI5WLJ1bgZXbMqMdAvO3ZWE
gbxvWQDrDbmIWRgfW2T7xW12tpytCkrySXnjeERkeEXo2zGKurlwTptqd/1h9HhJpVtiRvpybIHH
hy/BbDyU9nhCRgFNbHc6C/EIgvg0OlJ/tIx14TMhteMIStZG8SWcU+TFWdIEc9iAsHUtVLwZdwAX
Dy4706/3nNOEyfiiwzGDyNWPbT1F92WqONhvYTVMod7byA9Ia5zTLhTSugmDRaKpJEr/FwGmUAsl
muqUB7mfHKcpkeD2BRdY5qYBrH/iy+U2z4hShL2vPQ/E0s/w2rEc6uHZEnIeQZYA5sgCj/De/IQp
JxjPH5M4lhV5gO9vK014F+WUDsHeRzJgHayLIQOCOBQrbh4U2nnQiUrDEo8Qv5HL3naqsKaEpvpS
YR5J7qni6cxmdJiAbao9wyCHhq7LDvkdER48ptXHV5LzBlpNekUo37M9+UnCOsmUCTLovsLrRm88
VffmVfT7ArTXF3xGolwyWLPNP/WnyrbTPOYDpJX2c6FQgMBYQp5iqFDoAL6hFYl5HzTFq7qEs4HD
0Z91nLdrjOJoe4mLrkdXUvNplT+3Ld1VTSKpcDcmefmhCZdbhNFu/yquszJw4hA/dSOrZTkXySmo
wN5rvO5aUMh+aYX6QQ6o8BTIzW/tHf45EqcuE9P3JuDNqzbYJRpgg8GzkziNBBCcDoKR/ma6hCRo
8GDS9MoUIapeA/UqhXwY2m9zQbRqsSvpIhJmVJYr0gzCdKnAreuZCvLULAi1BGNikYi+jb9lJwro
lt+y1EK7DJIZ3ux4vSSXTxoEhNW/40VrE0KR5jrZxpQXBPVOO9JnZF/vtE3JQVNrJHDC2HzB7J+C
5+pqqgrqsdqY7v4AvX6luWV1WhaE2EbVJAoOgdeDjiBcM4M1lsvs/LCrv0SpLiC/rRtwRrwNecAr
kUcIssyShiQPDIjQyHfu8QH47rckdbAtqFo1p5EGAlV7oCfHBQJ+0K3bnWYBe1OkbiZSYvZbDelh
JiEwRoloMUIpmKzozIAnaBMo+UH2vQQzzJRaW6vulfrD3TBSAiTbET1/bbkbKnWaUEe7h1ogmfZT
gQNwaqXCXLu0RE6YYOUHTLWnCEmifqUmeeMsPsV1UgfTlUBgRespBdwK+X/Heh5mlhFqj8/FhHd+
m0fvKQvNjWZG45LF5UlcRI0kAdIKx39bCOvh9WsN+FHph/IUul5JwF7NO/UkQYF65ilJVbBy2qqS
9AWXXi5Pd4lga19qYE6jtFcBE7VcyjZblRFP8iN57rnj9FcZBilnXItxF7IUdc1r+K2aDdjDy0R9
v5sgSaNPZ7yOO+mwjeGZo5lxrHcgrB1Qc0Ju97Q0ZqYnx2N5jVhgwZLRdImNV8+xuBTuDLwHWA1l
h1qpC4WrW4TlnOLrx0DfDY8fOA5MLVyrzCXW8SkAPcJPRYzZBoSohhtR6s+eYVq9OMI3mLgcRv1P
NsmHZ3ZNAh0WOxJ56TIcERebm2e3s9xWvjy6MhVsoALoIsARj6kX2gxZ7ETbrZY/oLICjmf6hQ9c
/v2ytlnoc82fvsXOH0KlqWS+ooQhUxQzmth4/7sgI28F/ksSt3zLceghbkEx15y5n/MWaWlz3Pn/
QSDYbFwD34X0mw/s9EJiAUqwkqDsm73bK84CMUCu3u3V2TgWhVDPtFZ7afDTpVHA7xrArnZHO5WF
eOOjqeSh1dcgFr0/v79JqNP+iyKJy/WDyNLbOjzYaUJXX+1WIXOF3wCo9Yzs9J98vA3NS0b/1vJQ
4Rp1/tTQd7R/hNfYUoHwkSEpVykbktjs9jjDwf6y6G9CF1zPTwgS2uF/8Z5ls6qcpmA4Q51F8gRv
Q837RNwMwz0h4uiSCyUB4Ug2AT/6dTkYZJY9EFd31hWLjJ0128edGevvCdG2DOrZV+f0ZRUQOv11
E74eJXMWk7gKgGTlY3THSc2WyuzS3Asg7t1Qky81U9KHU4k6JeFgDo2X+5Cc+PSXXlLde3CS6jPi
LislXVM6MNAKmr7Y23cLMGiboIZFq7sZ2PbaOMEUkMUp9s7hbReQ8py6RfeyQNJNrMy+Lvy3Oy/h
YS8FZYDJXH3x2aWNi+OWz2XEtHYICBg7YJ9nWu5ky8j6CX6/Yvh55i9e5Qq1JawrmABXTlNT9ABx
kUkvnIKegGI/1QW5ftPKAhhfoo9RKdM14i7SuY+fQYqD6Nd1x0IWQrDwYGIIW+yNr38eSORGhmAS
V7cmVG1Mfh0h2R8Ri3pjbVqttuzTCMlUre4PjIQ20/OPw/xz60/3TVVaCU01j5F1qRLQcRxHKwAp
fLysVz9tE/U81d/O6nkRN6Ot23nNDwsc9zLlPBVSNKasjQs5gyMyZzm9/pon2333419PPUbSJV/m
HnGiVU6cIm+HTvXIiEqK6BEBB/Uwx/MYNV2TypV2CByk52Q3xwGkYx8Cqs7Ajsihrs/L+IxvDH+I
+mgnW/mMkEp+XRapkHByrFRtp81dGuOzmoLesxYr/VieyOPvNaJWh1hl8Uh3c9RbPnry623T5UqY
7SY39Cf40z4dCQQFIMbsH01cCtDV08U3XQoUO9e59+466v31q4GgGit6HTqBHJ/NtDSGA3jyAHyz
EJ4SCWpWtn8a/034lRmG/CE7sLssWI5U8ESHG6o6voGhfXMnDT+ray+P/YPM8W+lgU5jFE2qB4y7
a17PqjOIdy88vvGdND+63oVnx4hgiF53c2h8IrB4NlA384gGd0rS3qAgOtJGM9Dl3w0skfDZ+P69
KrrA5dPcy24Usn5Sb+P0+leFJWnM9w3QSz/qV761THQu6xNNbARgfaruJo+c14f2ojX7ECi4sXl3
72wpcFPg9zQulXHGsV4dFINBebXArIGm4K160c+9g3JhqddDnUXR9mZPnXHLIwyO/MeS01DDjGWk
n5rJy6s/lfFTLRYTJvQfKs5qafgTGVeF5V4hz4/+qpLKtkDuJhpm0H6DRBr3y6TnjydEjGRym6Zy
mTgJZNR/5a9Lsr0n0ImiMQwPvQpAb+kMdgS972siOfAyShM8kmLZuTZ4ZgYtM0Wuzw0Z7BGM8IaJ
6OzQZ/do1cRew6oYAS+2eVY/gTfxjXEPrtLxI4Ix0D10htGl63P53Hp651s41/1c9SNoWu1m2I1x
5BNGFM+0iLqvzgfldCiynV767wYaNAdSW5g8BzUkBiu0U9UtP35PKv/wiJH9oUSS+VY23TkxaUKV
lJ3f3xRXMnnIPk2PmFlA94zBLWZcCyvxXnQZKrTL1bT+MeF84tKixeRuxxSI/jQ/ouGGG7hJUn3n
VjxrNLboPxZXY9JDd1GNmLe0AaIlcvvLMqW2uODrvSsrUGdQ9kMano+2HmKRLPOFs/ToPHSvS3G0
EdV6gjnFCpQlHBSZJAIgUMkSSX13/FooPtA8ifjQky2/P0t6PMAAXj+vRA2gu6qLvOUDmEHBgI4r
s+/Tug9f5LRzIzeFK6e5Pe+J6z3IzoITKNlxSWnRQki+FSmNLDPBUuaFogn1BqAtUB8RoJhmZyhQ
ptqyVYYWocIvfoDJAW2d63M24WrU8HYjvycH5Cs3kuj9JeJPhQGFa3VRUAvEtIRlxAEDulodVntl
pbbJqmwjDLYkKfs56aZDwatX4tBBJoTAkn7tF/Sf+JXgBrDwc2P6tVqYdYdyy5xEeP/9eDCOb2Mt
pZQlvc8A1t6gAVow0DnAoZctpeBL3FCEhkm25LroxoBSf0L6pINGwpL/LqyAVchhK2RvmtDANnV8
b0q/pvZzRnSFVdzB+3guZUE/bZvZKoYWVY3aI3PFWBbUrjVoHqyJRXyOgNmwqGG3aMnmQKVZ2aSe
NXBqEwTkt5c7nnOgSbVAKV1z7pTOcEs27wYjI21kiluYnEeGahUzJXa1TaJsr4ipNb57lzlBGHTC
r8bSxDJOfivsec7tbHF6UYWwuUC0UXwpc4mol0pim4GwON4meXEYiNTeNmHDRfZKeKCHqef80tK1
WNCnSuOwc/4OzgigvQI+A0fKzlMAItLl0CwPazOtzbWeb+1dzeuei3XsWYcDNsVqa2yNCedpFSka
5Yccoc4hL62FySsDQlYfXM0I0o4jiAXih4VcnoVfvkdak5ulBTegewROaBRUpgqFRkt142MEe1fY
VYVaDsvPyHfL+WhvI8xlxSY2+lKrQ/k6LRrZCT8uIDkLqbC52cLOjjl7HT/oNUKFc/rI7fJGneWw
DAG/bsw5NhJ1fX0ewhTc81JNIdcdJQjYllSWQ/RLzAk+/YZor7R5igQaPrmQfBmDqmK8rXuhRxgo
+pF5GueqDGVFlLr9YQJZFMb6FzFJ1lJ3OdJet1ycu3z0OVG6W8xRirWciSXZoXkt/EvycS0l5oVe
MpXQXAMmvNhgKHxSV981LNqdiVxnJW8ZFAAuTpDUlAjkkTIF4f/XlvP0H4B2jpXubQjiCujPlGiu
jIAZWEhMFu1HvY2WI+oL6W5zJYFMzcrC1ACwiodKA+EIhImzk9P56Ai4LHZB3K9XXZiL0+bzkube
qoDKjfqmXozD4+kKoJAQ577d3eyJYXsJR2Q/CtOQOhoXaf05oF6ZO/HAB++sto7lwUGBH9bUkJl8
/jfmDVMcJoo2OSxUCqCtwK/NRKPhOsybgrvMO0WE/fFqjgih2GPJlMXfyy7Hh6CzkgBUFq9RtIIc
0CUoWL11skpTuq/0hcLR5j7R90rBplEOblxJ4DUnYc1UpFwa+mBVJo9rYdlnlYw24jmxUNfQPrh6
IOgCYb8B1yDjxwul6y0nDNvUQeI+Ah/o40+ppITEE34yi0bXVDgDyYq3oBTP27LAtqlvIiaEcAz1
cFZ54UT8MSt6y2ePKxeWWs6Zbmn7zd75q/4XHJEzNu/cdVMDJuPZPDiQzZA+cXSMq4HgNCkKQ7xB
hZ1fKKXXLwe3iOzZqHftrxkB1Un5E5lKO9vLC2CrJ7xyMbE09TaQBW8gnLgpJR1kcJ3rIvjIQXvG
sBJDr65me0x8MrsBFDOg6masDd2IBKLNpZKu1/ZDwpBqkNuHce5dEUwVmCEwZIXID9xUDf9IJ1/r
8W+VLPw7hy5vKXoUxJpONuShDSk5Q10Fs195IF9tF7jCxpesaC4TW1CHkjQUv+erg87sDQnsxvzR
pnvGNNGA1Sa9i3yIdsxH1lg9bokgYR0gjOaH54vy6u3IWmrBtGOz784ccUjSoMEsxvPwqq83QAhR
xV7xj9N0ts0hLh1m91/iSZTRTBfyCXhckbw+ysqX185XWqGZ5V3V/9/TiCPNiX6NKTo/a5EIeoye
M/S4/W1FeTYvx9kqO0eyiy6uj4NiMIunXlglVlla29hVlND12xY9YN/jSZnxRclhElWsxS7ZMW7Y
p+E4Do+Lzv9hG+M2qdWpXLg/v1r9GX3rpWit/93pAUOaR/my+mYWgC6OLIQdmwNI6+XnducOeUMs
rhJCdN00xMSSmM0+m9Axqacn+kIUIwJNSwdezy9UaBLMYKQYo+c4xCVB4IektxHFY3/z0czrLBOc
r7227dVNy/p/L/xEajjrjObsUIF7NzdWotzubafKD4jK9SP3mciH/JiqgN6tocGNNnwk3x62w73h
T2NAUJAhAP49/ns8qmTvYo5RdC0FHoCjw5sfLgJTk9JgoxvhIg+MkKVtSHtWEumrKu4R89BVlS4M
Rsdn5ISl0LSU7c9A6pyrKRwpTpdzcYeVrv4a32Vkqnro68+cZg/3xcDFOIweV1NrcdPVYKqaSwJH
t/7XjzlGhrvnFvJCSTyGe3NDM4n5UR/oNQ7ow2dWB48UUYVPqcDGWDzJ+v9nDRWWRaznvc4HSWiv
JbvCMJN8AvlUZ4owkxjOWOgY4eYYVdSwLr6rY1FvEa5oe0npbXratl4Rs5vsSlyAzAW4boDJN8k4
799F0ruihByNzzfrY3fsFjfgI04QBp45ZvFlVtKLl0nXV1SIWmGH6qMfEEt2RlvE46+lJDjtDkWW
yEX6ztGYpyed2T6nn0fMwHcmTBm29IHCHt2ziQ98//2ymvJK7I3PTR1pXs8B07WDJCf/bTqZCZBt
cqWKLW8h92xQGQVDvrhD/V2vTYtLKY5iRQXebYdgqYsA9gqGDe7X/UG520FIsPHTGcNQwRmUV4pL
eDPw2KMrw04tdsSiyIHye7Oh9vXAykPN5eG60VQEq8XPtAfQw7O2EbuJWxnG8tdWZT199CQMoNnf
JUruyOeYXUhu6JkHiuJNLSGo8cbGEPfh5FX5OLmigKdFKFJeOID2+YZHDCX027QlscRnq8ee4EV7
SpDIK/31yBt+0a+BpLKwEg1ea2dF+CTq8iycjrqfib22FZ1M7uDmyPFWcz5L3pRzH70vfhb35Vci
b+5M/jm5eTW6QL5ot1zX+keO3qAP7Q4DnqMzP4+d7xB3yh9sqxZDvwNuWNMPm63qTH7HEy3KMype
xGchgIvhUEsVdw1K/y5/MYgOqTpCTfLkSZnFhclYjF7z7pkWS6JrhSissMeiv0Girqy35yNoQOQe
HKOCPmyMrB/cqmI4rXBRdOF37HlZiNj1sgxa2y9bodFGbdgyZ/RnXjgjZrr81IFwet6Es1QJbQay
vHplvyivGtYlwc86jIbFpU8cKt52OxgsI1U+iuJtQCT+NlYKyalRRL40NCbGJn2VnGYnZ7HpBzP5
FGD8Lf0wNhbu1eIO8rMXu8AGet9JQI8Y+RvyXVPgKXCNgl2vegjkVJCtE8FMB8QJ7NQDAqfn4Mgn
Vp8yPWkPi70n1tlBD0hfYMqi3n0SVL9UGQGWt3VVVogGsIdy2QeqycCTzJftEXPhpe66T/jnegX5
Xpe7UTFxRp2e/RTwv5N0t2JEUEBWk0o1Nm+HrCxMf8ZEpRMWogdMQivzZZcKJkmv/1idYOSn0eGZ
oim6ePDT2tMExMcLbKV4V7uvh6QwdnmU9Eh2A2TbfDkxarsFRFLMJa84pEovKb72wTW6jpWIKu98
ieEUwMMelRFGXEFMrLxiUjwvmnG1wyWepUqpNTGot1veKWJ7Cvk3A/bhjWSGQnYqDFI/zJLuEkYL
df/jKukWNWQIB6zO4rYLBIExdaxI8qR7ljW6qnKFYl8/wjlSFoOp5dWiM0XlX7wLnf4BNHA9SYF6
l2oALWqueKlCwyzLmaRCr4rHxgTGZsCwsNb9GXK5uP5y+qbIG4PfxYFNYQPvPQJi5EYj8l1a+Lz1
ru/UcxaS8tXIOITVtBgc9Eug0we3RFifpfkNPi4RD5MVMLUeLWk8v3gGeMY2RXQ9Ir1+Kkdthd93
TipuoJhb63S/zZzkMcja9oldb2xUXGCfDv5wgHiD7JVtcD6+UbpQ45fM7OEl6wd+fZ0S+GZUNYjC
YleFWuGlF0nvzY2hqE9hrpjlIH/S2ltyS1zLu0gDFjgWjQ3HTbnBLqPpcWtJfhFvxraXwpc2LbP6
CVUqRN8Zl7+c+1VizmpDLsXLx0B7XCPRq6YFfn8Sx1m4jTkvaHAeZ6DzIt4MXiSM6bKs4MLebLnd
YXQteTEYxFvVH/rykYQj3suJEpOmHC160ZSNROxi7AIfUJ4Tb4mUkDRFgEODV0NnTbZK+1S3xWsf
hkjIL6O4aPS9C1QMIvRdW3Mdp2cotiVqMxWl7mOMrNYfcOGyr1SsK1Uh5+OiLfsQCOn2IeoCrXuD
7ynUHgyciRr6qp7GksAXHM77GjCRvGp8eLyFx2VqEqzkdFbh0aKG4jMneQvTRx51fIKMEmzCgUjT
z/+Cq6ylVg3nq8ytqDA2qC/f4VMyqsnHsMI9zSxCNJ/91OB6K4jqsYE8vxS8QHjOXmzx9scSKZLH
IQ+F2ku4OWn53n+B2U7y9MI4SGk2K+2mPdgCzWPet8XvxkJ7MErdrqIl8z4s1jaUb7YIRJ1RluXe
xR13eSTVXOC1UTTdi1HXK7vo/QZIZp88qj1T/8fUhfTxa82y/0f8AnpNkC4gAz1GOdXb1DGN0o+4
yoqx2cYey2qoW8SlO30zN6p5B5yNIuB9LBx/qMwHmOUq3Se1lfkeSd6eX41pYpIPtTgSjtGQFmJn
BDvrpbSCpOl+pSjEmllDVfUfmt3p1kEl/040ZCk/eYNmb1phck+BqvB8FYTuohtdGS8KsCAPaLpY
90L23XhxydU4FJXZgNMPbO+d2iMxCWvlxOAOtatWQQyd5DqSWlecTYQJZmhR17We8jxsZrRTGcA0
GMy5Cyexq1FZJCXhRenRVIJxOtcA4CPLt0oBstOe86JGpy8mvhGJHoTf4olqdp9WKRxTNEA6iwOQ
pIGLWE75+WcPSFSVYN2dPpojWwT4Qr+u9SU5olBOwuW3Ex5wtTfd03SpSeEb8qvX/REJsqXzgpGN
O8KrX8nqZDx/NnHvzLMACjCD9uCirS4xq+Q0IyurQhcCwF2F3GZQFGe/jfbv5dx4WnQ+BZjEmjvK
l0+f6BAoHS/88ZbzN8mUNUn/C1k8Tx+jNZ28tGSBb4TQ/I73FZx9kLylkbAS/MaZXjfFzZLt2D55
6gObP3Q/SEmnG7RcfWqJOTUQYI9UlXFwFspMzfymK3e5+qsYd1FIbzs7e7n2V7gE6ti7BFqwExYd
4ODgDSQznssGwmirZ2O/7KXUjD55/ANJVxJiT6+0NCLE1L9MskMxFS3XScfrv3bNEXHBQy6u/Xkt
RSbZXL/QT8ULpaureRmmQl6MH8JCXRPKXFLCyi2310vfGNE7BVX4olZUQjlNvLrDwnTDMssBFpcO
WnDHs8hE1+dIhT1fEppltX7Odu2hExXcH8BccWx5XgEjwaHD3UP0bawyB/uWSbG9/VJG/v0X+lZB
zX2BQuFM1Lys+IbBby4EbAMhQLKrHU1PduCKQQc852d1/VwwksSOfJJ/vklXQ2vk3+4Lw47GMrvN
y9BQqwH2zMt4YpbJAl2JwmlpPM/lOJlFL6rCB3STkQgenzXpg70brOfi2s4TchXUULZegFmcvg+E
0vwyVuyrNke+uDCUSUl3nv3UUyE+MVWodQkMtRCuPNUQYwOa8f0MpN4JvMZYEqtYdXEVKK1v8ofU
Gyzdtcs/cSu6TqGVdb71D2+o5kt0gKp3JIG8HmydPgSZoh/ZKaaxBE1eNQrK28GL77QMgRhYtOtZ
Mv8ttKBAY/kSJA3T3yfqajNy8Pb2TfwuZX8u96qcwmKWT+4hxN9XLJ0LWvh41bpFvfDyRYrRQ92E
Use2LLh/ZGtdgBYAnv1pxXFBLWdGpZ4aaM44oYDloIChPM4tcq3hQ2KkfomOXYqujWwpk23kEArr
jXRUOfU8L7vDuCw7OB2h1blDI7l2Wb0kMKyUKbGgemCuCCP6+uzDmmqX41+K1VYtFl3ysDfIIovM
JetWNGVczcxeE20Bb2S6uUFbGwi9p22pUEulfNqNshK2r6hklHgEznJYwqdVw5/YSxxNuxoqct7m
97X91ivRpT7rqH5FK/g/YGvDxmlMdmSmFn9U9Wi2T/zbm/17G9kAWxX55l+ExnjWysmu7NtZTmWc
9AGHorsMNnIFWeCI3knScfqxrU5keSjgSFHpnLCnbBkYo0scd8QrxwzbP2S2+zOCg0xEswZXfQsH
/F9kVMBq6bANaFD4eqVzwRvp+vKlm4Of7HU08EnE/6pE18z2VZAA3UbQnj+djf68dDsItZ4724fw
ZOWtkzyoZukyOToLsX9qpF6G3p9pEGHeXq4fPTrAX3wU0bV1sueyquYAPaR427CTdzPnHWEwyOSk
067Bb6+sg+BQVP6YNolsAw0DzGPIhP+Q+bB/bkeFn7ifqcbG52Oa7eTZqlDLI8N0AryEyBJzI+ab
U9bR1zSDPJCIBlTuMxH76VmGC7S7CAUByH8z21laYsUuuUCthYN1a5gasGuMXjctg3c64wDtWv0F
cuOnY52I7G/qEEARGq3kyT6pbyDx+3mo3307ntGq1U7cK6m3gOXt1wcUlb1Ywzu2Ogj7pfWYsvbO
uaVrrWMxW5UMaBV20a7yMWYli+Byo8vET++n3eVrz918EZzUQKrS2bClufZdfWlMpN+heBCqWT/b
7nmTmq3fczBg0p5fljq0pocs+u3m7BAAwxFirbUXdCeN/ppkCmgF+Z5krb0CVfLaDgXCE9+k8Ciz
duqR2+1kgr11Kt+aOzKHERpdkuaCIR+fNEVTIvGjEvFxeNn6rr/b/ExKUVIvbntKrh7ZiXIcMdLO
hFYdvST5sblMQBoIavgYOWNTrZ66/WEF3hHIYCOcxJN9E7E7N436OdN840ETf74oE/zP82aX8qc5
kPPOJ0y4Lsd0z+b9ODNiBCCsL34Z338840XBCG5XDu3Y3eb7u0gbpo05g2eng/u/7k1lB2HAx8HO
3KLV+ogZfC+pxrqU1x7Ot+1B6c1lLz/Ly38wX7PwPnnODvS3rzDMx7c1sanC2p8fzX3u/w8hI0+h
MRzazKQDFAhffHD374FNlElQU7eKRYatN6bD5EPP59EheqeBmv4cP7TtaSUtPbLvAuJ3+UxWn5zh
DUpXXTH/n+fQPDl/piyeseqti64vvi93EdMS7KL+FVR4plfTc7QDo9fujbL3EWEhgZCa/1hNLK3x
WR5WP0VnaHtmxDZsaALmeZIT690ceB/JRk/ZvKSawO2EOllLLDkhVe2nPqU0yeyiiiB9muYmDrxl
R1zCIMQqkp+MWR4JLoSa9fGCBww6YeBh9vRiLHfUc07U5UvRaUW5g3YhcE1i2L4rsvarcMt8A8PV
TWmiBrpTMC4mtFjJliIz4u+aRVPdHIA/yojBqze8u3IVxA0lAsJWho77e1KR8ObiqjvpT3nAkgbH
6moYZh9uyePe6gzf6scEVvZ/Qty+UBxAsNRY19TzNE7Wp4Mf/o0i44Qbuz/QVerUCSdbq99fM6Ds
TW+Qrj8evG6tGqYcgxsYz6AnFiczO/+wFZMB7wRxWQ9ZNao6vjDKIKQv6ggJwdPa9D5HaMUw1GQO
hSV776ktnAvszhYpf0dqixHEl6hjLXFps17JkGZrn38slKoUwGPO99UuYBizESTse43Cx+TQowXo
CBLjvsIua3N7cKDtxmByw4cGJn6psD0hEut12GEiKgFaFYZAndLoggi/tEZx0OHCmoiKpRsmWR/E
xEdDlFBuWKwA3YX+QCQ4Giup8X6B0rj2JAl3hNX2aZGyEcu4bvBSkoiB2sECFthlc1vq4g8M+SX5
hSB62iWpUivPcw4L3yXEg1SiciVofpq7js80KVh6hohWX2eRiQTKELFaZta5B17HdBEWeBtbngxT
mHKfiXSAoL4tB6Gz8dsscyM+gtPY5jSwSxa4Vfey1nd7FVNsVqMv2z163pI6tbY8I4RR8ngSnCLE
w1lOFx6eWYY04jIj/aQTqnGHYEZ8Es1ItZL96nkbd5E7b2yvIzK1AvHCPQLG1K7KZLROMvvagoA1
AlkBFKmd9v2vs4NC9RHDnB05KgafC4ZOB0/GC2avctjb0bbJWS2DaAjj11Rlf1iBx/tT6A3w5UCY
l14iva89rhROZFgvMsDvpph51lDJ2fDhhy+p6p4I1MLmf+13xDYRu0Ybhz5zAodTPFCtNBoHE4z2
wtJcl49wn16QIHtmES3B9fxtGKB921Z+XNoUhZ9fvmqGvt5+mDRq42WVzG6jOA372hVhIcsZNgok
W2UFIen9NEX9cqLRGt+pl0CAndOd9GYLRUuhAtiZJrfgdkT/kZ8soR3sf3zkIwLhE3df0XJ1N4Vp
uF0j+zwShSVoc43zXT55kODMoaHxdd4X9JFaeFjSj0mO7LjcMdmmAaD2l1q9QnxR9gbsyvHRcA67
6EqHZp8v7cvCIN+HJ/mYcO49TfNd6ImBTVeiWaAY+jPDHI4grGLXkg7yXiJwVfguu37lN3U6s8Wp
7yy2/NUfcgozu+XU3kFxnAVhmysrNqOPeleqt1+H2vuOHpghwC/22H2Nzu5E5L6m11AN0F6z6mu3
st8kZvxuXE466ipQnvuawJDKAS0a+we7nBnhuiRjKVB2ec4cVuzaTtxJF8sZF9p7yLMvP9r+FGTP
uJ+nCl1S55mAvpiS44tfnlSH6+iVPmb9iJn5Ds8DjOKw5ABoGNxzLytVmjmASL4fex7GiWEwB2cm
ZivLoWVodwNnO2SGLHClVume3q7AJjKBSgL9f0pQQ1rVFMDLp8MkoaQe8ioOPcpWw0syH7gUXgKB
SpfpyN+LGbYJltsCNQOOA9UssBKQJizVO7lt6z25A2XI2o1Y7qy7Pu35jQcs9F1Tuy6kDpgFCS5R
wDW9Lc9zdtlVl/4zNSA74hCgOgxPaU4qXiv68ddJHnrZluADcA4G6wX8zV1XyjyuFjkwkEMkpEaD
rBGVS1jxROzxVxt5W7HthUw8ltvtQtnregFhI9ld3ge/3H5+Z3nF0X7rJdOdqGoTt3Lh5DefiU51
TkwhlRtI+pUaa3UROETK+TDDv3hUyA0VlIApYtqccpgUm26oAdjuhe78gTiV0/KnmPG0jyPgE67Z
Gx81ibBLhghKBfefXT90O9vNQ3uxtkNH8BLOE9MW6m6r7Cqi27TLQPBgIF5AQEoIkEcDAmTFI7h6
rOCErEtR7T+A7yzL7khqErLUwW9BteUFdwtb8+L0ok2WKo9RaxG8PVziyHt4AqXoosl41dKDTF9H
Ct/N40+v3LkiwK4uQy6QugQwwqN18TT4cvROAa6QSJkRLV2C9Col+0bUgArB3VsVx83ow4LHZGIJ
y8qHUN03CLw91UdVo1jWGo6j7xaD3odTJk2XkJzs8ZWxlazczSDBLifI1kIsavorxdgY0I+hkNCL
Odpp00hTTAR3VZllgb0JUncRCOC6/yoeAvbNk/GYAhbY2BSDG6zk6PC3EN4E+0pZiqowRfIwX0m4
C/5HjxLXRPgvGU6SqBt8p8ABCXgNA1iURLCc7Zo86iq5VO64X+enVf07QmMMBLqs7g5IGCUjg6gP
t4vtTi56dy8nx3IP4p/JvJZJt9bLikyTKjgKFRA6PNkZMB0ly6DvcfE3ikEGsCE0PcsRF7l0Q89M
oqGkKwewftK/DKAWl5nKrLnT8vCFw6ftGi6tlrbyzxhDpjNchmpG1yDa4P6ezdNXiIGW9aBlyCn0
kApm5yht+Uy5avKTmdXnJBnJ+Z/Ylsb8lgJ6cWCvZws6QKDQ3D3J7VzJhmNZRmfAz4U26+0UGi4Y
/JseFDhKGC7e+gF9+0XQhW91yTM5u1E38/ty3ftmbU+m+6j6LkEPbuQ37aTwlh+xqYQ+3d60hRaj
HQxddMFwls3BnFzIrBjyoBfNpcDcJvXW2YDRIFC1IojPlOHIIXDUsgu0EJ/tvooM+H5Jrv1n4jRw
xkWTp1UjaBFg+jVOtkzhxB7KDcZNwMzgVciNQnr4kHsXnfGIwb1P2t4fPufgZxE2CHdagsImDdYd
Fci9pXPfvmo+BcrLcRqrMyW4HbxB7Gsedn/tHhmerVnLS4fvnJfmRi2J5ZJaWQ3KFLPClxDTFZka
SbltaKZV0IJYgITopotVz8zdPRvLWH4mWUYokd8N0HGbvJmJkbLnhm1GS6nyYkj0oZ0qEjo9uv7L
49VeZZok0EB1I74QaUtR7b80NzJpsl1a/r6oeEkkv+6d/WmfSvvgmexA8lF3TW6MYyyE3WdHcDcr
GBEGuHdyHdtTh8S7T4W4d+M27vDIOuMoghJM0qkyd91mW9y7VI7awekPzfKxFRuFVZnSh1w8Qvx+
HGT/GO/Kt1ONQmJ6AYRDavjqJ3SGdqR6ZyrIZJac50PCMu6tnnAeydT9+25IGK94oTotnoCcrsWU
JFSELmEkmLdpxJOSdwMR9MH9lIFc5Xz8C6FWIiz6bjBBAEQIXWiFGEl6/o9uiYwWVhoGQj+EApRU
cIrrn87pTqmjBnmrXF8JEqmkpRkw2r8+x6W8hzI4BJaJCVGpneGkF8hdEwvJkuEbPG5NMCc8kiVs
GU74bDOBHi+f+2l72Idugcl2WD0tcdAv8PLJTMvIOK3Q83NiyUi+Kd3zbI5Jf4zyviElCcCZHtw6
tmI+0EuXwIenCqaqz9y6EfemRBcJ4Rbs4s9ucK33GGuJJNDe8Hw9vhp5ovrjbD82QTJGz0JjSfT1
0vK8pGRAcI5pE2gNF1qM7Q0IRn2KIKT8lfmZYlZkuJPQ3kzPsXCACnBIKgZiWjWeAQ+TnrvXX1OO
PRBQBwGG5k4XHwaqdK152nhTqKXLKmqUsDUtiH7QcMhqCPvnRmro2+SVWJS0CHyr6wqbNqhKt6/N
jZRnO+ZgGOXEzclOIR+zlfNHbhD9JHUWHKKFtFxtWINgKVJerq5UpIgVgkEL5oOyjqCHzqpna1mm
WmD3Xe03ngbSLpSF4tVeVKbAaxndKjL1Gb5a5/Wnw86NKkaIbyC0djHRqu1CBSAnaMYRE5k+nzuu
Jw1UmVCStJokgEuElxiu7dJ9mlzR1CI3qfzC971Qrn6MGTfcscDgkRrIeRETHLFqf0EqJM2no+zj
QqUYuv+hu24WHorcw9M4FnJl3QFIi5M3YImeqQAZJKbxUWY3nvAEwafWF8zK6A7EBcBVaMtC6RZu
wm8hqfu5ShmlumG2EBt+iP0YWicfisbGOGUnG3MEZCTRMkaf4MIpsUFTgLFRRbtqRzH0+YslyIAx
vJpOn6305srvaHQxHlvSjzSP9ZZS93o8NhNUg3hgvyt63moKly1Gj+7sIytqqeXkGO3JjAlV6de1
UPzKagg8lNSQHm5EkIgw3TKEmWGrhHMSit09obppQOx+bBXZdRPk+2IiU1MMrHmH/ouEb1PkRRxi
jG0mDO8QzK3FBA+dhedtvjzMEF7+Fp3ZvABNbtBL+TNAMJkukRpC5mPAy//o8QYzqtkJoTQE4eCG
Z6EURf25z66VdTEM5XMPlwQeLgQTtxhr3BQ9vkYgzH3yGtac+k/bF7/Hocnskt0TyRetdqG5KofY
6k2feYnGpsf5+0Nguk/ptXU8BLsYd+Iek1VGs1hGnhFAHcR0YrAiL/7HSFD/E0NTRUYr53bQYT3D
yswe74w50/05oQFF5UzhmYOYAWPFXL/yomStY3IVy9G9qsO+nEQ3BpNxYnPCfFlyHkK+WBXG19Gl
0HLW2rtzgd8NJWGexUp0vIbC8cDqPAQeEBHm4KpPiDZUzszIAYT16UbEPJM+M2YyqeyWf03EdrzX
zrCVKhRasPYPWEXVrT02a86abOqtpHsernaYdIszoTOcTXWskGH8DFtTdLIfZQO1T70vs2ITAxXV
J24bNZEs0VnpflntAKYqGc6fJuWcCwkTF+lv4Lu2EePxoFbgIZ3TRnqwroJWFXIaLy2JJ3OsPAdW
CCkvZBhltfiLisZ3j9qYQ2ev0axUlzngmuhgNH5cVo526DxuzvU5hhiQQXpsLr8Cx1UfEFJKWjka
1rIqublEliyIc8in+cgx5vlceQZSaGeUvxaFTvEPfnkuZm4LIZjfntRa6aPVhN/I9nt6a8FfJFnC
s7NQRpDmFsmUduByFc1exQj7TyeXARiR2dNwB+aN37HHPGiujN2gc5Jqpl02u/BaF7582R9LmQy4
V03wa5H1Tn5JCNZtdgdZW+cxvX7/s0fzaNHrL65OQFgnq2OXB33AhSfQNkTmfYPOxgAbvOx0Iico
MbZuf+GJ//UXsDEr82GZ8fShaERvY6+14mnwcvvIKwOS+je4V9zcxTvV5/c4/oQ7mdv3N/wwvXVG
uky0LtAVEF9wT1jkh7O5Z/dKpv34G0yrt386T9AHw5tzLr6Ag03XLnoupuKzvIych5VgMqSX7zGL
Ig5vseDJhnO4P4ag1jRrmfc1dTzr452nLaYuMu4TJP7qbtLHmDuDZHWoP7ljGIKyjhxo7Cnga0e6
TJA66llp0GlzTykSnPpE894ggOYNT0IIfPSSK447Q7XA2CLbKj/3YYQdL5xjS/QRT1s4jPIKkk4d
LiLuz8T/S79joh40CYH0Zp3+GVeJjP+xt6zt20pwxKUn7WOGHWD0EOIITe4R4BINYnQVN6I+M5Lj
VHnw/qOdf1A65ht7cB7ciixTd3jNVIoEhLOfFBazIlYYxBxa0EV8SC6d5+9X0ZZWPz+7SGqlJoT4
fsmvpStSMo3DwEV3P3fwqX/+QTEMuzSW8ZUjL0IJoDLpk+Gt3IMqe5j54bQdsKMNd6JlQlOIJTyk
YhVnUEq/vha9v0itaqM6MqtfBDf7mOA/iwJCtOOyJs2uS7owuQfZDIG85dlxgc/+SN4uN37VZ0sO
p33Rn4FNpNeZKufa6IbG8FD2W/zmPpvuuidRcGGbNiY6JSqcefVx0q0C3sZodPNQScUigS6HkhGk
7kI4ZtJx6S9fiaPP5G9TK7bihKbDaAdDfJNvnn9+TG925Dsi+DWY823BRLqM4rWfJfTq1+eC9ax8
uD+5qdta+V5QRTi0pVuYeunss7dJxhDIeBpAfsEtQkRH3yMcjBrVB57u2j5CsSPEVn8yFTxohxuL
40vH+R4Hlg1tzInKXSHQp+z/gZ6rTpIzZf3CvCwQPyHexhQJsGGfxYEJAfbjqX3qIKVUUkkJQwQC
fIU5Ysp4or0M5edCW4PMBTc43cibT0gRd55+eZDNZAmQIl5BjcUQcNABDxotIUZwTyG9Arlr+0YQ
DHsv05e/mRFJUSHNtr/I1Q1g8XrBKkPI6H9KRMiPfjGkVR5FVQhOvCxcsruji3wsr72wCH4mvRW8
Xql+ws6V/YxWAu4NhtajNcnhj5bCEe7jB5hUootnKz1w9XkZg6JCYqgEQO1NL9V7MIT3tZEAkEUE
wFLDgwuGewez8RYxv1dZafMclaL1ng+GELwkQk2afHcVOML7JhgrUz8n2n/xHfm3X5WRdmhwNrhm
xS1HGSR9vHYsn2QWcQbryA4mipGoy1Wug8m2/VDJYCRbcsFEg61R3U6So0gx+g+7hYcOyMNIhHgz
3nGszeksC4A90lxmo0OGvR1jwDNEnIcUkY+pnZIN+U6Flb+7V5T5RY0dh67c1+24APs4v1Cqkh45
42L/T2J+NlJzAan7CQ1DEa69iNMErOCRVBPJL8gRfZTSOrOokmwO9aOzpATtTZJG6WR72uIaPwbb
MXEogMGHoOlNRFlPBgxfpNuKJ+ymMli8o5Y2MkBJTxmcFqSMtM0iLYLwGp4A3ga1x0bgR75QKzNl
cKyzrIJ/BHSnTsB5CpNirLcGdtJYHvt7KkvQ0lVeDSbNq3p2LX+vyyBotT6DUaEGP+SqQaV5kYWc
av3ICd1FqH3Vj/JrOqOI/WBqSUnoKOXgowqOF9EXjl92Cn2PGj6vEDNGpfAIlSVG6yVs2zKZ3kfH
GubmL3n/NlmpgmSxRL6Whn64R8juztMo8EJZ3j30ORNkOVG5FNgspLOM5gsdFptGb7ob/x1qx7pb
HROiX72zHYyhZOdXnbPEvH9MZC+RBntW79q6Z+j0g0aDC7QuFaVX/NMtB5U9Q0AeyS922tQuAQsb
TerkoHgcs0i0wNl3a25cFv42BU0iYdqPvxMHnNKt8xmXxs3hCACMTXzKt1q2+Sk7vyJNGESjtkcF
Qfa3c0/4Vkkmfj/Pf3oJB1aTpX+N6QUUqU8BQITacspaH5Zrl1JuxHULy5/1rqdMq11qcQfBM+np
eVB1EIOipQ9VOCTk6jjiG1IVfDuqCXvdL8yExAMIb4c6xDbHgqN2cyEirG/pHnJdMSULiHJ+7PZG
oP/ZefyMckh+nX+iTIUfxxGUGAU1q5YGut14Cgzz0aJp5tG7NY7SW/4P+mRksDTq1XE2pPULSzej
LnFieIDOJijiXdlSnB6wPXcGVtCjRBdljars7ouPX+aI8JMS9maaxSvbsu2UneDRwOCZAUxNMsBd
0gtlIrXrsq0V+NHvKrlUUGmfGmMQK/KIFg5bD/NS00ocM30X695OD5NsqRLDwtWIYI1xe7zqD+sB
GxjFgZTYx//vew6FokYV9qCXL9ykRKXCM47ABbVo8/SFUJCctQ/AY6lI42sHK47wVZ7mAcJy5hIS
y4LcNMhHVuLTjoXkOC6aPiWy48OlsQ6IFB6vcsjdAg6gXTt0Di2tXhINre3WK4lRghaeKyihoC8D
aJqWtUn42PkYvUAeH6Wg7ID0TnKfjCHwHnOMB4ojiwIijm9nKiE1LN2Ekkpt+D3p2DJ/ZcITLT8l
2XRE41sLpNLdhfI1HcRZWBN/4jOn70rM+IB5BrtBtdBcsJvHmGjpiB/Jrtv5z228cHpeAyqpd92c
B6kqd7p2KtHywDT5pzNLH5DSQfVW1RQw7ZlkUH8Uvz/JD19/rTgaHmJMnQxo4LjDHlxgbT6PEKfC
WqHBKvCS1BgWfY/Rck0WbzyjTJwNuwAcDo/O7cbN1Q7sXiGjRR2Whx1TqTMzZAyHakzSwnMPJl2z
uXxys3YsZRE67fvWat8RQ1hUVOeCtUna4slZm7pJJKc+wErWjdGtVSCbIrDhMOSHH2yIO3TWy9yr
xKOqilKsfuT+AV75X2liMlXLNnSOXsnWAbbCwWj3F71d4/ci8m2+oQazrxMqPk+9lUiQU2r2yGuK
WRKKPwTwdu0eo8oRucQp+xwNsEJyrA94lLsicTBVO/FcVfAZZGip5CNm4s9d+vRF99T4vWuYUnt7
RjgD66pVGbMhXaGwymgMmHj8oSUbduWkw3tUteGwrFSKCAWW3R6jgFIAS5YfeBkY4i0mY+Sk9Y/0
k6msV/4fHbqIXKsqJxjO5L//3/q79Eokri1oTQ76CN5rQ/tnbGs6ijp/Sl1TeeY7auJ0CVhMAN2z
LLFAemC0roK8PztroDYN26UbmR1X+qcXcptE2sQciWf/gE3cqG3aeBR1QK6L9ww7UboOra1QcPW2
zlpmqn4KWwh78ORSUw69GyO2nhX9IusiGVN4G/MvXmsblGIq8Ml1B2Iv4uo548a7bOVWGQYd5MSg
HA1vCqD4bkEkZoWj7V5dprsuhmofeOAShP95cNSRk/yfZ+GBqAg5l6F+Pk7JcTqy2s/QZULiQkT0
vOiBS9d0eISINIBWuHVSSA5qC83Pyq7AjlT/2kzi7Qg+RfGLlhPMoeNxY4lEXrNNkYxzHiW6a8uG
2ieRlGDS5r08vzx6r134kp9650/Py6/8AbykjW5URRZ3rr0l6Mpz6zsBiZ7qBdThYpxGYq90MyJ1
7Q/eajX3ondh7qt8Wi6Ba0ZM6nsOpLy54K+/kTSujtm+oo/Q+uBw3tqhpgHoLr/C6JNplJDT5cLS
ZnqVkM0XeIQA/B8umY0Gd+5uDxC0D2aLteiSEQXsVP/KIRYSElfIrcjLYc1iH77Jg5ia9ihSgD53
Db0X6xXN8lSIEuHtzxUQak0WhPDJHcYzmawBYaLbSoM8D4IvLj3tjFjFk+xE3iH/vVMeUH+K46Cy
BZ4mMcrDkPDFZFrXNhzXU8NqR6dV7IFKvb60mWgjxvTo8Hhsq3boBO3Pr8fHfikSyUZECZ7ej+/k
XOqfFN28YSYXB5m9sKWpU0LfEUj/cQakJDIY1zJpfSimWDccVk4F3QDNFu+G4fRxu+CsHo2bAg9M
oWFzmxZiAWfSshYH5KFLrYKcgFtjK6qiKO/yXO6J4V/1ymQXTTZ2y3AdFw3C2wNBrodTX+HsFxe0
sjHQzyJCehGcmB131v8sF0J2V6dzr7EbkU9GSJBt8o8+uBeO3pBGVnaU0pJwnIYAddD1Ns3TNk93
ALpwWmv2SmHxRbCOtSU44lUSA/DiGbFzWoWFKf6wVBfqQax58o/+wj69s4kHtK1xLdsIDEjk6/wP
b8ErFgWzwRHdZWyrzmRQ0nby5Hi7t9X25ebuhgHxdp/yUwo6JA18VWjBWBotZyNrB1SHNHzhcHnY
5V5+cfWtDTVhKpKcHZUTMmUZfdNN2eMnM0AV+B/tgWxaDpX4oHy8X5bNBBgMK68KSOJ+1ehX1Pq7
1Qum1ZgCgcFNja62ycb6uaMdvDGWnitxtCt1i7vFuScndZ+4yUYJyv2Xqaetol39xJgF59NYRL5P
1fz/mgi/yxc96IRqRMr+DyIo/3hn74+TwXzV2EXoZ0YNrAKIUA2mN2wjEp2nelGIJ5gdT0jKNvnL
TjDnkglW9rY4QqJR0VZ0y2U4mWOsfZVO3z5AUcPVLpFFJPcWG4FCnvF/d3BKfcB3+WLh0BMausww
bBVzZQabUxMwWNt7AsTWJQTtpG9Y8zWtQrfJXQz/O2eKLDirUTP6I8kZ4ojNBatC3y9s5abB/vX4
7Gk3UbMIna4i2Xvkx9zsrCALA2pi1euC6DfoxqgM+G6N5itFUpKjSMrhvomqN4TEH4a3VDL+qNqn
EWKqiv+cKwOj7kywRNemMW4acG9qo9axWa7ONaugiXe+Ub9r+Iw7cjmso5htYUkjylJdX8v79h9X
pVqSUVQYVlMzc0ceig+7iw+I2/kpH4FHDoVSGkwO8tBmEGL8xVMhPjvtEyFro8SXNkkTUBjtY+2p
CrUD9DMloO49FkhoqXN5TSXmNB8JfE+KjHp8JApLyQto7BP7CrRZN9uVpMqsPmH+ZQfBm9YdzYa2
VhRMjWoJe0bTdMj1iIqWQiZA3iKSlOICOhSeVoLw+DXKg59dJwnE1dcqZ50tNgj1eR02jsumyQNk
a3IAB1PnQUcwDvBAUDPz8Nxzm84dxgf910dFRby47onN1bx89C6y32NoCY+d2BG3PDMLUwghZvYR
mH0KbFiMk0GIENKDP6gOiiDWYJH7DAH/IGsqd2IL8l3XK7PZOfB7hkeckQUp2j2ks/G7XQOHu3+d
3uC2bxYxWrA07KtNHKfJV0XWnuAsTBig5kyvzu2YriuUP3sGTnDP3bimGdiylAZk4d9ryjweVySw
vAcuPlNz0UI3K8NnQP/q9CSMBTItWOrNhl5zHXxVpFAgt1/JhcMZjyLiY1OuyS3cabxihNH8KJZx
kzedVf50eglKIfHt2JTVb3CkvBW2/eGF1Fx3f2LkEmr/f/trXinc2YVn/LRA0ptS9jJW6/F57sE8
wESSRHRejqVn573UEvEoxW8xum3ucmuOCBGd/OZngC5UfoYRyjU+RmZB5ce1eM5UBJl6qsCtvbul
Ps2mvxn+aSr/dIQZbKA0TKee+tSIV4Dqu4jGWQieSPivUb2Qb+jzELUog5Tpg7AzB4KoVXIZKJC4
VFTOIHG9DkESQoSohYmBPiZwV6Jfb3pC+Ib4lwfXL60N7a+8n/EviuYzyoLtLELmTPP2qnqV9jnT
Md6hdrDAmCTX4mL+yCOwhCUmzjBqEKQTIpIJ8Q1+LzAcnHwgOZxMQND70MSCxo8oFXSJz0dAtd22
3NoiEfA8ME0ZIsYVr3GfQUO+DyfI8mLb//gxepMiab8mJEcLFR63SBeEk9YWlBk0MzhPJ8ABOOF0
cE9qyrumg7bv0xX6K+Q8UqGW2eZrIJfD8D9+H17K39KHJZZ81w8ysVhXZzzui9xsgdjJvvoYRGVH
RuKi6JruTZrc56MgLhyQKekjMgehKn4mjTZCNCOKW7ZLA1YhrOISpN/c+OATi+1w9fEPFq1ymxuT
5VHwp8qlSlvZOCa9xxhhg4O1PlgtllatJGkDuTaYq+VQGQtvOyZM1WCNqjJxO4jFy/dII12Gg9Q1
o7ydHVWG/9955qmZw9EqabQ8WnXQySD0ACBj2XTBIjwOcl02oIKUqCRQjexBIEetDjKMIT1x8wkk
gvsBIdxqUBZciU/P+j9cTu5Zzj6aunwpkaSx6HcSBoENY9TnQ2JGflStm4EPkWEL7yvjEd9F7XMP
wU2+CuIK6Oq4Z2jT6LfVja8jOe5rueDgs+htAXGcofZlD9j8+izO0rN8QrJF65SskQDUQuwaK0pc
atfSjXB2fi5JRFxPZmM3eJazbL6kejwvKdjnkjokk0jU2sZk3UPGeA0gSeZG9H2bg5jcmh5OjjoY
8sWktKjVBkSsfqQ/XBYPzkxfUc5+KsMUGY3GOJz7tNYWQGJwXokb1LeKiPZVA2vE7FrxhvfX01C2
CMRm06w1tPwiUWUwVG6OiWPrJLt7yG9tPa3+A5ggFEpM+SbLzYY6D2x5Q4pct4Inf72zAfTasln+
k4xPgDF0oSC5wIIlspm2hRBdSqn1wNdd3SPBasS1e166CcQGwgYYIvkPe1Nv600XehQTFOCq1cdq
C84B8HNkx1GS/3buBN9s/hXgtb85zIIkINuSRv3W7/ICWI+M8xcjjzzNUyjDfAg84M8fqhAEzG+o
uMQulBb/+ChRs8dDNZUALXoLtXmNFEz+5or+4ewjMWtcduFtqfzmWoPKD9C3fQBjA8gW0MXq3Tv9
Li19e2bePY+lhF/Vue8+HKNuVZX6pP8C0K7IAA7J6Iv17IgG/T0uVpcjb5HV88VXMf8N75kesJJM
B7WQB1RObSSALpDkX1irTwADRSDKx97W5Pd71wXGcCXWzJiNQEgLsCrbgKqjCSYaU/iC4L1noT2K
akIXvyT6qxs4/LF3UUhczlUxlVS+6j3lTTsYycVn1ZYELt2p3BKQi2DtB1qsZGpWz9gnLkwtUshV
OSLM7U1nb2y9DT5t6H7T+hIq5RwVTngmUKnBx9yKoCKJ4iRaID0TVOyedwoEggGtpFhjWa9k02x0
j7RFwfsggwGqkU2a/RRg9Oe4glaqfEqznO+IzMC4zKFc2qvQiMyzo7zEQhoU8ksFWCgUHGvjsLNC
e9/Dwz/7QCvN7DFeNAOIJgFBfrgsSkv6XumL+2QQStGPTbCqXKRNllGCVJ5rju2mESCphcdf/vDO
Zw3InERr2Te9QzfnVGv/nfudkZWqsbclqiAvqu+IO0oxMByUirtVVCkX8qY0jb0EPHcvshCGyR1v
woTYBcL9RhjtS8KxFTjvut94dgUNP71TisTTPi2UApCgzn8kwIHZYTjp/ea7DpGPaoToihGN0IxE
XuKWVX2edgBWhdIx5lCw/72W0Oc43L9fDXGa2dvmMJV6GSX6RnF3kiH+as6yfscwYPjLxe2T/hJA
RVKAI7oc7VP7cZWe8pGZBdsoHs2vGep/zKcFL3xpkmJY5VaIb7AYBuObf9LHgnOd26FESviC8fGd
kcKxYKiL/mZj0XTTZK6jD83Pie7CjVPdgPBIBhJDHrIDYBp2oy50T/z17VHvUJGB9uf8Jnuyb2jh
+h2JW56snV0JtLYvUo7O2uyLEPxMTRT5i8uK8q214TYI1Fe7RF7PERD+kOZD+QL1gbLvdKPgyVx+
uY1NjkrjXBoAlt0ULJMcZoXVeiFOxbNXuPjpjKqd2hVmApttATKVQi+srOJ0qnYSDWkrZBhEnRF0
atx70ERg77HSrGPIgflDY9L9D3lHbvOWE9+axppA7MQqEdidtcKYBRxJqiefkLsrVCzyuuq4GxMo
RqcmjBqeWGghtVpOIGFDXBIAqRlyK5e8ZfefoiM6JTseNmehv/4JCu0ivcMxdV4mGBf75/geOWdN
1eJr2hnkHQXvUJiMNJ200VcjwImAhciG57ECYC6baDcven7tRyS+q0WsCXwjdcpWBUZahnEdn9/G
YIcVb4z3N+jNVXQ3ZQ3KRQEOaTj5cDew4Shg3Lh25bRC3QuJ+ugoXfq1TETgW0p5+tLlrBxvHxcZ
yp7YV4RAp6sVhjFM9XSOOyoYK/PC7/2Lj+bplqdVsgAuc2LZpsRTaUXJMhS0xAzX2kD8fEvk/0xk
S9WbgW6YUuauYff2kbVb1iQ3z+Tiokum4RVfUL+m6Q3r7o4zbH5HLO4I/F5aBYa3sZ6bMptfuW9h
tvSm7KF0XwnT3/KgNZW7gJuR/eaD4X1esvbj6nXx0/PxAKTNUhkIe5k92AxcDxpiDnUxoAVZZEQu
z3xaGYVG+xs02M6Hm1QWp3sbHd+jGnEujDRzAITRBCKp4dGO24HEmr1ruleVlp5V4wrTBUkCymmd
8JCIFfWBfhp+gPJWwJFojeUJWh+r6wib3TAQxTGiKpEepHXhxelefGoceb3AIz0MGCHvm/Pgcrxr
3cgwlrKS2U8PJE1kYRz2z4DF1VN95Ppa6qBM3NGXFvnKZ3wksKF7UGFE4bzcwqqJGjKObnev11A3
Fm9vzkWIzcUBg/HJ6K3IfRORHh4+Hp28jB+rAaDKoURYlXZIKnTne8N4VwfvEt0yBQLc+h5LtvqC
U8FlHZZq3r9eE8attmXIoC2Z8jdG8u+eK2QuVMhB+qMKtpd0uEFlGW5UWcdVq82DT2QrPNsCfMfF
HXzCeFp2CywVvT13E7J3UMSG7nhPDznYVq5tfh9gPI/2B76kB0e5tyX+AW/Nb3Nd3S8nwhFQQ7o/
lCnPXmqyk+dnu6eXMexY4dtJb3zKq/T6hEddxKpVOVmxfk+JQjh/DDoJzWRljWj9acCbUnF6/ajs
hyVoLcG5Azsw3+bZTWWxbcEWoImFhEnjkndB7J6xCNiVqhGos2kv8B0oFJZF5B6Fdqvpj0WHkJ6z
748jerg1O7xtTkYcijm5RD7aDUKuAxMyG/tETUFvUv+sqGvwexXOZybsdBaDUYIqVgABR/iDKv4r
/xjV1RxXgQjcvo5g3pCP4WhlrIuZn8lifLtNZBa9O/MTou6741ljKIaQERJi6F/QL9UxM1OqI6q2
PYyaT4bZa3fdpGE+EuUvTtvp6pf8UgBczRdkH6wqE/uZSA3KZsVrud+MKdtXHXKVnAKvlNZkjBRn
/FKpEo5tua5M/CHDUCPCP7V/U9bIwei+xQNHGtyK3XFLS1+riGvOUeS0DErz32X531UC5Xl/aG83
jrkavJhtrB61tHkwVrRvcuRg5jn+0aCU4kD4bd4AnKSV7xGCDeiu69qHPvtyqao9hAhrYbFYWMno
XznIRdH/bm+p8XCj0bJqSx1Ri2+QHQXjRlsxmvfxZfQVMIeTC5pPb0v2OesnKUfK/iIkRLmEZk/8
syh9cJR+26TFeW+DMwOxwJkrB0zQijTEMDDVEKAuWdY6U7L7nn9jn3pSHpwu2a5q1AUSTpfyISI+
p2VK5FWl6toILr8Zopxwwx/ct2DEYiITWQ3xjojIbwjKtQ0pWqV3ODvfkEdPAnZIac/H497eTthD
pyychZP6t6/VxI5bOEXDs7/u0oxPHzj8RKfDFPzz93WNK/QLebZSzgbnIRGTDoA4k/85JFiQ/U9w
RjEpk7pctQei2eNIGcYnhWzbjsKEnfqSb96hC8c2in/XPFSxEK3qiuRnIF8ok8IFiov6dIsBHgfj
LMevEI4wOwsbD/zVJZqiL/BtASgmiZ1TYu5AS5d/LkPx7qg6y1d668btuf7QZxMDUpxzjCQ86Eu4
Z5UdGa4AtsAg9MxepqtR+pr1E7mYKLgNJE2u8qah5I1b/EKCSQe27aUa4rEbTDZ884VoHQefXA6f
E/IBvWWsFZrEmttwwc9V4nzq2oLUz3pDS4nhRzJzdUTD6j7WFr65JyR5E+z1S9t89vanVfzlnU3R
tTEWC3kw632m1DWuqIlaBDXjbbexRhjvCIjujK0FPb0G4mTHMe4p7lh5v9jfr1i9df+YS65Bcomt
nuXbsKhd+6ezJGeyxof4Rfa8L4i3ZiW4DMFe4yDXBQZAYYLtgpJRDItjFiYZ+1qKH7cq7PSaqbfY
gOnC8c6g0aMPKnFHv0wJ7YO2slAItvAsW6S+k0g77aDu2QPTiEHaAX4fAvfPQSXlQba2QhDL1Ei2
gXxKRVrTazv6V3qEgWluET4JVPCvsZ75YqtOYARAvhQ7bYnD7UfWVhgAZukzY9VX4q6kNoC5vFoe
t0HWiNlZ3ujibxebRC9BWpi8Q62saZtJXoqM0bYguw1Vla8DWPX39s0MuNPY3hctDQ/nwMg2zYCI
q0FrNZoBruc3c5JZaVkPjkKtkRUevsEfJtghp+kKXF0Wf+PcOnNcIGuHPPXSu0Qjzbr0wHGs+5Lk
JvILJ3xGPd+6D80L3Ek78S68mEhLpFLJJFiAwtrtdQsFBFUc2DpnmAHigfuO/mXn6L+t6hKgrRQz
dhgUQu28z8vmhCEO5FdItoy46Nq5t6bpgeGE1bmwxijFUh2c6fVIbrmV2TXy/I06k88Y7+fiAeiE
xmKrcxqnCvCSNeVnm8bLaq+janxny6aLr3aN2HwzkQzx2RwbEe5blHT2iAN9HHETjCqo7ZnvXFj1
1zIBgTK47f7+xVCi+PuUo/dmNqX4HQSvOk9B8BrBn+79+Lxp1JJrSFi7MmNowXwN3l8BTopf7gUh
zGO+471QFeRIZRUr+m/9+8+HVwiSQe4MXP8dcHInhdxqT/WGlEC4XYdGNrlVva72Us7YOSXt1T/O
sXYK/ltKtppdVrKmv0YGAbSAOk3WI/ePEC2AZStkvgHkN06EoT0PLIF08p2UiljwXg8neMO5xXa1
mbuokaRWLU8/DqHEHXQNho8ZQkF7Kb028N7UtQ1yobP45GtxUpXL9QBL9tgs7Ch/8Mo2vJUaGL51
Jx5x+/aI87y42U+Zi1x9x1GtbAGgXgevD3g+vlt9RU5DjpjRD3ky0H4PPX68lr2HdVS6eHosujMr
9mKbAAsQ+neyzwRSQB9nYOUXiQY6u/Q+1V6NHOFOpdvIJAsyLNLkRmqqDWdHjZaIMoFb+dxJ/GVs
45kNUKxiZ3IsR5epHd9S7PRL2YmZpl+Nw9i1TtDZLUjHObFPN31dOw+oGM+EgcpT15zIGwNnvdfT
754Hvf3K76l3SEkTN75m8C68HjrBKjRVA22A2R/uut7n0AghuSUSPp+kjMVuwWL4H3wbvGyW+Ma7
yLdSzrNZrdiE4+e4SmWFikQ9lGw+D22NtKdZuihx8ow0Y6MgXG8TAWKH2WWDAq5VKkeRwVvoLDu9
1zz9FBjermw83B9o8PgQsR8r3hatslrgwLWl+RZXgQbOgE2V5n6H7r4ePKdyMV1aTgQgt+kJDxT5
8yCjh8neIUm28Pe+XIO1HYz2Sh/o1S1wB2V67aDim4iMbzQEz2w3KdJDCfX8YIx+hHECbe/wZwYW
Z4CiZ/rKCdlSrtskef8roxiiPREnmfeLrzCvwWk2sknjTApGtV/Hf1vyWDbdWVDKvfdvMgEQd23H
ks4bxKZGc5AL+F9gXu0xMsBgtTVFux5UmA89F1xrJfeN58bCztiqeFihVHDa1d3VN/nmnI6T+CO0
YIjlyGAGA1b9fQhIRz2y/4iLhknzkOSjREFcIb4cqGkPDExI+nqNzEIUw0J8FdR92Ef+uuF2/z/q
Tw2r6pzbY1cYVhJFXPgR2oaIzV9zRF4qZ3UkheUUH8Y9szCQJy4DG6RjYbssi3Q2TB49tXJfONmG
mUDewr4ULyyoSCIwZizYyOaHHWFsE7w8bv4aj3MRDhPzG9lkBDUT74SKHAwnEX3y/zsiP4PPzbRp
gyh7TwnNBGkyQ4JTyRHcvz43Yb3WdGnSslQUxSkmQASP/r/iD9/TBklOmrb4t3bDiB5U6peKmoUp
y55HvHF1L5oInGqdRVOqotZeUg7Z38ZiViSYfvKh38WjeF+yYg1P+mbHZRMRJHMudef13jphviQq
hYJ21M2GqRsRqMRLqGBjQ5e5hEyiz79rcMyLPm/HNAiCdv4iOlPOZzO2qHHIGTDE0ul7/iF1dIB+
KchLlfu5sMv+oaOEqgKBz6ze5Ak8WlR9EwITFH6IpomjaQenM2akuufWtpF8QHpw6hcV4LlvBtp+
KhOGYJaDzDLyeGCndteiGc2KrFnQQ0PkRCSSWsKNqAfPOI+kLzY2WUfyhd8J1hA3818EM7k8P/Ja
P8VL9N/4LzTb/5nzqjNcRPwVSmOqoqn26FF824Sk6f/sJ6fKHRCTSaOpd0kzFgXE844MkL3OtbIs
sKBJ+Onsrltspl/Tmb0dQ5cqALfp9S0jlOwALJGR2Yl1Vr0q9M6Krk5BlHqUB/pP5/VRSWJ61R1e
4NEbHWjwAvi3TMB4coCa054NnhVS0AdzA/i5Yh43RrnrIbHg3IzlVk4F8L8VRh4tz+trm6RD5Bd0
2pK28sDN2gD0Z7YFjcvIOKPHgx7JCqTWYv6WfucYlDgdaxfpzISvH8LaxoxTmsHSPsn1napESwhL
K4izmQKSFED0FVJWmfFaH6qT9tkulOnlNbZR56zm4qVOB/CX1hyaJlN3P4fKvwiDsx/N1TPwIptK
5yCBaPVxzjktdZfzj9dw6gbhCD6CIDpI7PWhJxoexgVQToigiRD5O8UZ4EiTwIjZFjaE+YVzGcPh
GNZHr+OBqsxwStD6al70CC1W2ulp2HZ6J84+QQr8DJEF8gzix2bYYFxbSYrR7ISmCoLzu2hsPWxX
XeTAMnlTtFzON4X0XNqO3xN5JJpT+b82jeO1buhUAW7tz2zpFDvsIKNkKeWgYbiEnPiHpeKjcDbK
IuKMCq78fBWyLbZsjke0ArjjwTUMcSMMDmJpTVqi9CKuz9Kfu3Vc9peTc6VkCAeB8fxlQTZtqDNd
RPdj32iLVC0GUWGg+DlNPjPeHifXcFbE6h5Y0yBEjcCb6h7/QejOM+Ex+OJy4PAAx1Dxz1FPCdYX
tqyYzZiK8WlkU/tMHViBcA3JqIxcvtjeaMbPC0as4EDbRSxI94KFsepXnJVWyopOtXVUpgkUeSWF
0cyzAVLCfH0t19VfAGnw/6t0ptFUxrrnXYKj5bB6xidD90zPRV+y6g/PX3RxzWqrl9w24XZlbRYn
s+GCZhQthO0wLYMLoUnlH3JB4O8Udp9DmNh8XyMSR6sN+wydb3xb9Gm4DvbqHMRwV3hzgLetxRaf
MV56W2jT6KbwzEYExCohwOJ6Ujn92ierePakufdkCpXVRB4x5jU131syP38dZpSpD2uyzPPsJFzY
eXNi9CSfpSpUmxxDk59VpLtkmyVAmHxen5FuAJlFCd4xGRCubskRQFcmIGbaqz69hQ7KZnkL7SBj
oBRYROF9nz7LFtJiBZvQMsT9DxyrpEoDrSMdonvDeG0RIzIq7VppX6Z6UcHWkqkMsfwE6r7R5SIA
NgCSBb/m4HTtM8c+YZz811EzLILBHZ3svDJQUdLggiIYDbJVc8sZHWy8Bc1duZoJl8wGO+3VJmHh
HiF6PxjkGDlwegWGNXBJNm7xvTyaJlxsRLq86pnXqeinIyMDDPB5moHeS1Kx4lyPPlLbFIERL4pe
TTV4Lm0FgD10aE3qxeao7hbaG66sqW5cDvAApD7SNWdJvrbUqRnKRDx1TmwN9Kp3AapHSMkdJJfk
TpBbAwXAQApSRT8SkQNHWZkxYqAAIS4q95liMKt/Bb4Veuv8aY4kCg0hCnBloVMuN79D0P7YuQLl
pLuK5yMlo59MVZHYSXCDCTwIXIctjKueUP1QC0L5rdYiYrv9uVYRyJRWmXONukjgx0PN/X2tmAck
ZYxZXqt4rQUBsPuONiWnmgpZ8Yk8TV1ZJ/hRrGa+OPYE6rvaYDpdk861n6oFqZHtLvSeJMxoUU1A
YEcIZPoDHdrUJfT5izTGUhRm/mzgDbMxXxcUhNUhHyGNVLY0UqSAITi16bYp9m+djBSYqfp8sr/d
DRMRNZa2rpxr4LGB/Ki+D8nemgJXb1hCkqIJ+nMf3OJoCwgYIh3E+Dnw80VVJrEOzoehuhE3joc/
AdQGFV6Z9t7I1cY4ay1TsOhKpX70CZpNBlYiflmF49SB7eyYSIfv8S0OrUlYIamsNOlXz84idxmJ
sF3nTSp24wzNMRNdfTI8gM+k1TAGnIudDxHjK5laIwbqSReuZNxhQORH7KZObWEHFRZ9PvDvg+5e
13rEiDzJBEPleSBNZZggsjHEGYlxe20NwTmXH8aJ6wktLULwSlylGpNUomm9wP8yJbDQ+andrtAs
WbOxskyKg4bVfV3wQl+P15ej1C6gDhSXJ/ehBRsNOTOk5k5FpjIVYyNYUqQ892+SIil93JEG0Qsk
bo7i8CRqbhsgaPgrjZ6puG/MnsdQ23JPZ2gU/UprHafQIMcJdlz/4+2Fd+r2UV1jOckOgF9x/az3
fbUXnLcMU4QWfHHAiawaSRDkpp0RpMxwHpQQsx88ztxoeAPDFXmb591WYhMd6zYH7gPStuganUGh
Ttzw/TDze086iuz2U8yrMp6IBXM7xIeeyTqeYmIAdsxYY6OQqbw5OMBK8N0AtXnoNanGnQRSxz9T
ju7RnvMKmQEHJvpMFw3ElIuWxlMvJfLCFYJT1Ieu4AE47nB9qenIjUp9mNnDC1wi6YPFTCnAfl28
hPg+79rG0gBIl8XYV9eIk89fLYiSECOHLrkDWm5El2yMtFTaTqIFAvIUSPtC69iHYqUrgsWtCsC3
DWLMPeNbKfzFEIt4I0t/duMaB/CEtGp/vUjwBF7EzfX3VGHjoGg0vh5j0KlQds/w9shUsoWSXd5X
A3KaOJ++XtmauDlBrxL+khtkThEkNk/SeaZuZjBiHmNaC171i/e609mSyT9ADEuABn3mJeC9xjH7
QtfRnRppFDnwKVL0gAzoPBiXa1MN5zVRjrpxvuWWlCtmv3IiKCt8qi9zKfY3oRAgg23xcf1xn+YA
3+p8qE4uMtyG4wTqeO1tSJ20Pv548qM1U4FLcAyYWvVlPAPoPDung4+qRnD6YmfX9WyYJ6oWOF7y
fT4QTYzqWZO+AEVFqqZ5mV46oMYzbSHTCuJzOwxmWP2DgiOmoUZkvU2RyimM4Q3qsaiYItk7vEp+
Ipw6iFfyHmem1fcURFt6YwDI7kM/pM2UCfXyzx+FU/CKPhg/t+Pv8OpwI1L8NnJSE1hjvPK116LW
isFxgdge7nb3PTO9IkaU/uhLyg81UgbF52Ho+HGbY47GYzuagV+4RiI4KWCzmETAUt1aJK/kzIKg
vizwRI4oh77eVPIwgYJbToK6GmdjppHTEVY1vMJeBiplUJyjLLz1WPuUyY/2FBaPMjwX2c3y8Qfd
0Ls4oPVjZ93EJJZXH+lnfdpWJgCLHiFmCpMRgkYRnVU+5pvKQUiwwDFvFZcqF1wLD6oM5+nNnYNS
JisKNxDUYbvhyY5yoHoWCQ9NTPndeVTLvLkuLRwB0xC11tKIkod+/EAX7kw+BkAlb72ag5xe9YtE
J8BaBPT4c+3pRwlMk4j6ELrXE2lE2udBAbFvnoppxFw88JCUE5Y0uZQNwzOfEuYWCN1nkqrMApzX
8MrcqiKqBxmxUdNi51M0IdQaU62nmaWHlUeb+i4VqpUMWusxGt1P4XSZmyc/gY2HG80layFiKRY3
DffU7RNotj1ojW0k0c93JbVNUlIn/b/xZhfsikWESzSgj+4xIZVp2JD4S9wnRmU2iKF02DeE3cy1
04xBnVdl2eaD4wyKknKg1E5OpFmy92Y9hoURELpHWHw4Fam2f0wi8JuGkjGr5/FdPHeicvP8Whcz
OLLUE/Qqaua5lz1XcQjdNMXh9ZECGm1iQhQHuzCMf5VUa2Syq06If1WExXsMr2pEA2Q0mfTZwBr2
sJbm6yCsOoW15G94oE94MIynKHdK/0qtMvc5t4sGzMryEBHqO05VfQahN5EU+yTloFBUL2CRiUp9
GQGxGmuxP3CoWLepEvjATOhciffTlV+7ZybJfy3bpjYfSJ4f7eXegk9D75F8l8+mBPBeWo/x161q
3d4wOolDrABz/JN//o8qGBAVPwrLU0sc7Zurm52fIJCYaAnZGWW1dvj7iD1QKfgLwlSGqTCMdEvi
DElo6ugfRgMoj9zHl/6C0lZBfLgUS5KhUC0VDckYgxUfSQruAioALh6oDMgU0OtBL10vvW0DMyKi
KcjM5ckMyoe7jHqEFLkiAj3hKjdL9qZFczY6+uVuNiCGunp+c1rv6kxZmnO7B/zW6KMBz/IKQYOI
WD3KrjJNetUsMQObujqjSdxjbjJbFIRDu4vZafSxR56LkQdyx2LaPbFhlGJjqZU7y9EwRk+4oHr4
bJjByg8Erox5xMj61D84Ppg9rpmgMWe49/jbBYKjXJ74/mzq9zoQJbvmNkLnle0Ne9hHChRRKUg8
txir4VuKpndaeUhsN+/6pJcj+tQzvFCft5llVAfEPw9tSxBJ7iUnSsjpJS9KaQyrGg7uUvjKMITe
5oaLbSXNbGmI9gu75beM+mnl7tQV4w7C6CzeOiwMjdFi5mo76npF7U3rLqsAQQXZblu5xcqURXcE
PjEzLzzjIvZ7unbL4jrTkpTiMqEe10lpbHblBcn92k/uCqUi+WznTKxd1HBMfwoD8bS/GEOOFStj
TFqKwG0pNyhy8nEAbD51kMf5G1XEUEMTL31z1Zft0G/TW/MJQVt2hbHUReyw9bv67JUQiHfJnBa3
V5GxQWQNXlq/X2TFSK1KbM1pq5ccqjcyhJLKrEBScDrQqzaRuTNTP278G3izGavK+R5XHKzw/QHi
lFrFyQsmVmQhSevKyz8PLQCXkkEr1dIn7rnn4xJoAe/S9MOp03qAtqRr6RpfpaUGyaR5s36geS5L
+50QUgkzRp1GlpoXYJkCyWqeJrCbVEbgyz920vPg/O9rbjlSRZAEppHZWzI565c1936aFIPPrbF6
DSFRcc9JbXLw+y+9kpyPTK6HsY1sRQS1aHxMla1f4yWJHjeLaaDEcjzxsPLnhpihLrYZE/SspKIV
d0V1xn7vlNXr3P8QebDvq/ivay1HMqcXWXu0TPb1Ep8+lSgmpm6w2QQkJ7v1qyZ7nwd/c81O6oPo
Vbcl9kAVrfJxodmyXVgeLYzcBhjiT3Ged4cgdt9oOyAFzWTT3F3PYAyaJAZfDNXqAAccmuNoMssk
KXhEJcEb7ANavYubHrkiHE9LZp6tP6AlKGTLgc46ip1Ecg5+0KDpRIaiJBH7IEiNQoWVZ92SapqM
g8LIg0yNqIia32NYfAZB+6iDCEjDiLfUhOXU6eM6VpJEFxjATAUUW22AIWL1SNoeoSjxJBrrCVqV
gBT4bfZR0iPZoK3jyx9DzYhFslxtbQZxqjIpQLsdtv8QANp+4r6BgmpnBO3eUO1O8p8PWRFmQB9k
F3boO6TpA/hpIpps1+QzbbzTUTWKCs7ezsRazn0h7EXDDafQJGDV0mlrIMAm6aWpg/E3TzjmVT74
6hRU7orTdujLXPfWmuNdVOB58/avoKGeSep3eeDBMjLUTYb1auj4arVtCKI/NVukW+5/JLgWsR8f
Uj8WzRAX6XHG50r6gKMF67a3NKtwtV9v/tsTvCO4hnSHCPR/9/nQMg5A7yGv1/IzWKQYEukiolbt
GWcYKloU8sCHjn9OexkxMvwvdvixk2IWAutzG8p9cPY0DXfbZtOnIxBTlWv4EFzzdm3BsnP5UHCA
9X2WwRaVhMEuf6RJ5lFcMdE/RRfuGRT+vPGbRDTUw3PVBTR0vlmOKai6YJ5ggkosfHpyS4Mdm1fD
Y6/2hur3hLSfxURltx6qNAkXeCxAfAfYtkBeAtQvQ922DiakmfzzqTGhmMzQliIrfy6ii+d0qIoT
bwzO+FXadLzIuyoE+CALthQ42LfzWazA/dPzQZRP/cSOVkkXdTHUcj5loVXXiAKTpNJx6Mgrpg7l
ZmQUrEoBuKMNnNoqxBAIirZk21s6gFY6XcAQ45inJrphdet1/r8xfNxcJoskcgeRS3h1IowLmpTv
CkTh/hT8WRixFYhyLeCDr05QBsgIbJOXWM6ClGKLER1g4N/pAsI0V8Ou5ZE5W0mxjiMrCOmQUpWf
gVd0dLeuE/l2jcJdQ3XNCAMd2M6T8Wux5Khrs0bohwwXNj+HQIMfGV0TclHjheUKbZ3i+O4EBnli
mgXgo7ErjKe5wnyO+RNcziTYSir2f3eJR2dXVyEPbqaFXZJjAHggj8fHwvQZ5KA3pamkRRspxZGO
VBw1ZMZrYQcBXJihv1COAa0zNmwPUsvmTQaaUZiew2ZradN27UKkXwsCSqcuONh9ojvZ1XmHf9Rp
kok/u2U8gV+nP+xW/JAm6JR1FAD6eMfMe5vLJyxjiTP/HZ2B1ojvqJYLgaL3lQxx50W4Ebp3s+4U
DWmKvXd0nKi7tnxGTfWx20EQbr5MtVKZ+v9XDoWCG4hf50KjAKz47/fm0t8P1wAH10VuhKQZVAEA
zxmRBhU9AVqghrjOGIEI2p4AYd9aanVw9CObLIJ5e1Q2+fPmtM8s+ek9T2fnTpNV+jQkVzqAJriR
aw0Ph0+cC8W1+GX9dPDBNbncSbCQvJZQLPPe9ZP6iL/D9dXCVt/b8vsiz+0qBSv8//+/l4YbkEev
GBll4+mxnAK8pdcGctgen/kyPDAnus6RKjHAv28GU8VNt2xmpbRXrSK9Qz/wChSSksoaFFSvFgih
F0aPYxWUNRHljwgJ7HKm35tbaMtKl1sS/AJL2NXsXPqcZ8QAkbM6m087Y0jQ/kdDBo77OtkabdkU
zUCinYSimgRkbKruZfCloIfQsSBxWntptIeae8fbiL9/8wbfBKxDiKOYfPf7h6YAEKfoDu+SdcQN
TqUZUSHdiQ1OCiHBp00/e7vkEPgTuYZt95gcbhUz3/2rnzbyeTWB9SNL1iF+K55ozmWPUvQa4P6m
zNijduUUXaPaPla6XccOZ2wjUyP69n8Mn8QwJjH+m+iiRwtSm5pFCLKqjqRRcikBE2IuSRF9ULWx
fIpYLWU2VPkZbvC/usLj+gwQ4uYeaTS02hupthPzB3h3m/xhZ0a1cO1L39cAL1cmafmqAYmby3CK
5rRvced5N6KRVm3R0e5kdHOL4E30Ff+hJMhtBGJTZyCfl2KZ8gx3EZIOw0Ie6K+D4Bi1u0xvyLtr
TYhW60HWZWH9DvlBoi72IQDBzOoQ/qrl/eWljVF4+2/3xVBFKg9lit3VenPuyuKQ2pP0Y+N5twfP
wpTPqZfXtpPN2LC6O8ge8OEhQ+qqHVBh2AuBFl5GKA8Z3CRyYUwVCXwzuR/c5fbRo0xyL9PfRyZe
mb/yaW5I/rbe/pZvty55aEPmNd86Ry+SzS7BfPcCDcn0hAZiZ1siQwM7lpWJKj4FEkPrOUhkwIo9
HAAkZKgKbjXS6LnRrdPs6JCK9zDSFjcRvBpYLL1Cwcc+DCoKKbzrLhmsy0+4HtShrH1uV3mVqGsY
YQeNCEGnlZOgSKuBAxBBtFvERI3CKae9GARu26zbuRyWwhtjjVlSvIawpN5gbdWka34lz1tyPUJN
IE1lMvGo0i63p5lUxIUF8EZLH7O7csz3OSmOG2apO7pnMfkYbPYqvbli8j0xbMbdr+/URB5zepwn
QY3PK4AJqrJT9BqFR8l+xy2NP5eQ89oFR87GHtj2OSXynSgYmafQLj8i72COjXqMMTAmWKdOStoh
EolzaWiLtM3eftcM22DSJGeVD04d1ybhvtVQoPeDvtnKNaOKP5b6WyOe7YmbxLMUsF0uwjZXBkLo
/Rg1+nMl0wkBXnGlx1DyApiKaeb/1fYiMIE6nM+AZrdzfNqHTtajCRd68BFGFVrAho2MY5scbe+7
qpsZPqesOquWFexE8SbsOfsjBBRpU78iQVmdPcXA6Zq+CecX588UAp9EMMYqPAqAVXkWg9CYwyzY
0WOGsHGLoNFi1O7MbTFoPwIWL/g659xD14fOj7iGIlJURca6ywVgghPzON94IwUk6ZNTy7bIdMtl
4Kn7ZyZdg2blLIc1ibhrKZQNYZIbJSurFX6PlNcK/B3oSfvLIoHRukM5wUtmwtzezxbCX4tK2Hb7
A4P7LlT6aLbQvhTIu84vmWW/lhpVqNtBx/zoKTlD1uG+6VcCmFGr6RLb7omWogWw8nCqiYkXyQKf
URLKkQcrPBCx14VXxzG96iDJMiPurED+b46Ej2m3GyITUWDk7Bj8B3p7KFQRW6r26e1m/qAwdoxY
Eip1viFu3Z7um/hNbA39CHbYi/XXn6ma+7rE5TI1zmiAWm9NqSZsvPrARP2DhnED+QhJ7fD3hcP1
cBsgKpnOnpQp1lNVuDuEYHi9IvGHhCC8niFPehpLxy886ayq0GAOuEU9TixH5/MiyPt7J06/2oLf
90vaxG8WFT7DUvc01Xbvfp2abTW8UW1Xakn/49ItE4rDOwdlAO2J+5WySjVq0Mtntmkr9W880qhW
KIPW+JX+V5rFqmF7m0Z7Bz2hF+kb0ffgcvqGwcb/cNLXad9mY+H5wQmDL2pX3StfhWSt0fg3qzwt
Idqq7PKB7DeQm9P34a4a2IVEQ0B5EDbgtZoQtvHadaPme0b5d4WdQMWsD7duNvueGFH/x/TKSWqg
UzYyIfbOtvnN703myAjfORD8qUAXUzLW+Dgv0NfgwOmxnnOGQOX8ZK4vek2OZB3gynPnluJnMsLq
mnjxWZRa9Yn0AnD5WA0+16l33KgwQkE4lM6sziUSZuwDBY2aLsmEh4Hdw+s3o41SD1VXj3gAluQi
97F4q5UF/jaEF0i1mQ5fb3uIBErwX+Pw/BpxLsdSG+1Dg2AJouJ+dS+BUDqFs5xrs3gNi03bK321
55gxP6z1UjIkoBqQcoJUhARrS6iHNc63e59Im5yS/3onav4qdxFNQZNd63Lq5OlVx1irGTx02+sY
OW/7pF3SXHSPjuAJ5gs+c9SOHLxR9GMicKa+3h1ss5kUv0acM/CUe+Zs71tYS8gllreRsmo0whfF
U051lhlGfO3fBfnGttBOuDOGhWZNu3W238f9bE3Tow5JEWLToTHD7gG2bMdvl9X1gaLpOS3F1cYz
O66LgUGDPs9ecrlRliMvgzWqFTf7//5iCC6SgO09fzzwRxgsbORBXTLUjwYEDcqHGZLksgeEqBP+
4TngHGt0b1RRl39WndiTWAiRqyQhFP0zwOYcrBBkSwLuz09aJBjNayOsLr7lOUzkrHKvWtu6Q2/d
PDtx/28kwpolGjrL+i8D7kkIvPzMyDC25Wmhsu1YsrtSvpDVuvG3GxzwnSpjdy6wntTSqU2Ebgtf
Lln+deR03DCB8mMFV3wyJDXxecLr8gWsQ41l5HbElJfInphw2Y5aFo/tmc5GqhP9o4ByuT+IzENO
9BgwEIC2UtT42XXAyY8RDWjtLRStVPHC1SeoksIZhNZXCThGZ3V9JvyN1SKE8x4cCw9kMv+0Jqe1
oZBWq7Y/aYF3dhhDlimKvgkpFwqGbt32bzGjM03JmiB43DAcIBcVQKayae4oqCX8HHNDNa+7DNo8
kE1VfsXl4Gucf2O64FKFljWQc8648LkPAA3+eo0iznU0QvuImjprkUes47SdRIqvUAZMQObyiZJV
vyVQzLYZFTx0uLWukmtWoBqxtOzrWSTiIT7oyp9Y374zsVqcsU5eqLgPJUeoLd0QUyTtvIRSye9D
pO6ODg6gww68QhcXYe+s9FPkGjiqPuI64ymeCw7dhCUBSRHcY7dd+DMTPzBY8eSTLqm0UzztQ7lZ
5s15g/ZaZM8Z2EfAF2qEcCyCntsOo0txmb6JMW+5EQBgf4Ccp/5S4launmGQyppbMTxICgQ0WyQ0
X+einiMZch5qTgQ9/AkyowfxUuBrpXgm9fW+MTWKnOKkMXH8iUXyAt5LE6ckiSoK4KoJ3ywIieok
d6ywlohiHYY5a7K/aGrx6/hSRYmwl7Ac9V/Hg5SDsZWbD+ChpSllfN72nME8P2CwQo6E62XGF7ML
vdGpCe0hHKkodF1ALPEimUQ4uPWfbO8SiuiO7NP5q7SaL6/zT+JMjwA8TvUlKUCWZ31USxuVd1jz
9rqewdgY/7ErjSi7Oq70EcOk+i2EOmKKh7S+7bcQMrVHFtaI1LW0AtAJ1qxLJKTZlrLRvuRvCbnY
oR1GhEjjWYWMDViZEGNxD8QZ3X+N3ns+PHUw0e8epmn3rQacdjxwJTBbA2KVxPvjQP8c23Ylbycj
ps6/KPf9WG65PEdM3G+D4TxlHuuworej1ItoC6xl3SCE5syZpIKrzn6PrfWafQYmeaaxxNbNf5xz
7o0gUWGRNpQPRYtHrFj+gqEzc+KC8fS/SUMNCz4lik+EKR6+wVgxz7jcLNR7k6LYxrBQ3jralEGe
6NNUIS7sBQcRoSGCJzoXr1i3nuvObAZm2Ylq0M5CVUTCW6+aed7Cw6JgF5iM/Bg3uvEqT/kM6lxG
ggke5YBTJ+095aJZEEhL89k7lC59MviN2my+Ixa0hUVHOi8qGNddn8KKEvTEFg4GdJDWCoSTK9j+
sNRKz8FGj3Ve9hIV2hx20rM9LhkkToX5n3QRKEmT2rgBC2u6v5UtuzPx3lBXTy+aLSMQTSVk8Ewr
q/KRVzCjkLC5ruGgYaTIWsxfoQU8GjLNjKvXGYPHkqrkCsHpHivMX225uoNAWabeGhNWY94nZdB0
S9/9Rnct1YvQfDiuBYrTeDemxtcTO2fprr8vEKZmh25+m6If4FMdDa7uxRGtkLODOCb+uOrwVtwJ
IeFV1ztgf8217ebCgaCo0PuLX/vx6ilTPDLM5U216c3tIuwzK8hz6PuvULUmkxNXlBoRRmi2yUy5
GfED/vWfRmzV6NepzNOrLmC8Tpnv5LEXBkqgyY8Zy3+b0NAxRPmI/dv8RithHI1DiNfh43Vwor9X
xJlyYW9wIIPCyEAWINpZqwJ1vjoTAZt/tzx0PX7WBmNCE4QBaefYcpES5Tv7ZspQ3bhdlNhuhwXo
V+0vnaZrv2i1vIP7rI9OMr8FG0TzjyqiZzMz/eZes5nbr4QFnBZ2z6YngEq0VVMI+D7U+dISUiND
kFG2s1vzVqvyAB6xAz1smNvFYT6+FvM4wuB29uxU/W+BJDV+aq7fJJc7h8YVE7dc7GB7Kgtmfqkz
JNtg8rNihXY0qzxmxtHXxDijdL/SOJuLKVjINL8j8bRLLAI2pJkrV6YDLcXHJJWfkunl4i1wtkJe
7jgKyyWN/um7ZB7YzpbYhcnMGQNNfCwxMWmR0v9LZRDGc67ainPqV2owvim63sDhifYdhHmfA76M
iVpulBCMZag3PseS+joZEyXwuqQM1NMJNDQgIaHkYiKD3k6Dyd1vQXenPz1EDKDOuRxujCW3oguS
yx73N43+cIaWVLw0Gk1IObbLQCiL3/e4AXLCet8ZzxhhkO9IaQN5+QndrVZ3W4wauVm0alcdT45t
P+pCe3ciuZq7MO6fFegVKIheVXaZ7smUFdmGOLzuCczG9rGjt5/ARX551yA/8rjYBtkgRZmGj/IP
9NIsJPbPTCHBYodLthvZRzrNwwGDrjlVIfUhmOU5THf9+yG/iTJC6tINpGfe48qrxvSyMNPeY5Ls
cP5Y/AXggxduFOLldWtzd/rAG+BLZT1lNYOUmlO2eR3MMdSbFaWT8+ilH0uu+sDqzfKjzW/XnBRx
XLwWOaWtyEo3wjGgQojqrDFZcWfW8VePHOl9qRvyY+n3MANKhsrqeL4Kp+KZ75Asj+c1N1zI18z9
15M+8zj1arIef0dNtMMGTv/yBOUmEcN6psnbJ/aZTFkUA7vUG2t32iodFgw/Po6trqwP14I7n8gP
v4wEux6NmC414X+CWpoX67znQjxg6aRXU0xiMgyxtzKLdu3SUZwwur+W/FWfFxJIu9KYDVrkqdqp
itST4z9CFPt6ie1KKmJIOirs5BL2j+fUokkYPasrvDabO7Fnw/mm4Cz0c23/pxYJYsajevPsNnTD
DiZzcjYdOWsacP2xiJydWbAJSuFhYCm00NM1e3NO0jRTVJyiyoR3NOZVRtv0wygO6OFCCQtFen+0
0Q8k5k+V44yQanyRCm/P3W0k8JAM2WxK878PyCYZkNOYn89SlSsJ1YGAPafLzNd19Rz4Li6zWIcg
ZwqwQ+jENZX0CNoiMaBRM91Nl5W7LlRwwYrNcILzP/jiqrkEB3mCwOHFCnVAUZjasyO10dnfXc2M
vBAR0fjhNXSt3jxhJTQ1XN+VRyB2Zxdq+Bf32ZU5bVTVWttyL6oD5+czMjWmTTOatMFSkFJV7x2u
BWvM9EB3cGLMQGSnG6+De/q/pNtXQW6V9UNF1VEjNaOIfcvQv4rLXtVthsR1S6bAeZ/+l/O+lOQv
U8H6ViDJ2wJCrznKAgSvSLvkfLrAic7C1V6XYyAKA9hpOnKWM3vk05A/lKVAUyeuva7JWCpyNDHg
hPJ/XJXYmbHEZlnUm8xexNvmvzRHOnyN65g0d9bGNn3fbSFDhz4MDk7qQebusG/n1d1lCPU3WK19
pxZPKfVdt+goBjc/lHf4y1tufqeTs+WdKprHAfh8Vgt+NRVGiw44UOTLFwdjKXeHKGzVBtrfsReG
tYmS0RZGiNW8bChA+N1vVfcCyOdYgbHDTkup+xBqfDWLH7ex+jQebqBCAUTvppTJGwrmuGDwe6wu
72fR1xThO4EEGpB4RDFMr42XY1tTWSBRYj5yaXyM3N8unrFu49nx+mVuXZuY+LSQ/ZwkFMjF8hY/
tf/gpBzAiIyHqx5IisbbTPckdKxyH7o45uljux74JAdVch89mEy5fn5sAHAWLpSeaZRdo6RAzwuh
0lSx0GmcjdEFo2ldQlopxX86B48pLZ3KhTpFZT79VR2cQ1DU5qh1NLB/qIXZGEKxuasvZ3rzDFIS
Se8wh8iuOgflZMEzpDztRNNWmfW4mClS1VMNHTgLdxGkHf4NEveuywp6tiS+DdG3ctDhfnccHjuw
y4wBMewPZqW7kayZgE5JcsdWTQPshPY5NVLp2njoxDeNplGWwU2MAclL/V3nfL7CZ3DciVHNBLFa
VLJ/4fizYpTIDuSATQ396vmwYvZdu0urqnqjuuZkNO4kytlO7lbVg39SQmwElpxdh8QbPzJqnjPs
uxxeX7I8oVwvkdEMB1/ZaxjBXsopiiB8j8sQWepz9G22tdZ4mqs6S76BjV6gtcrnSUmopFq9JIcP
qVpyE3ioeVeGJUeOGOo0iHAcIS0xuXfvdhQPruPpE9GOXDvVWYnbim65xKw/Utvhv7+xLm9FCSHN
1FbIFN7xs5I4A49VHE/2wIC97vKxsUHLL/E3ciuwPNULgdI5CF/gaUILPxDnAN7lDIs+lPPoFocS
PRikTsHNqcRlzKS70G5eSCu+EvX3Wab0JTWJiNE/rCtN824WFL+XVvYAmC/2VAIa9SUykBA0+g23
OlXZsqO+K1rTWpD/EZylmven3oTXOcpCrkcYKoj8ohSikThUnQWOa4qusF+VgM2ehapGPpDBS/Eq
p2nlWIBOSzLOBAQ5fyiUDu4l55aSigGyUybkBCGCC/+iK5vFoTFoW+okC7tRN6WsF6yEFqU6iSjw
f0Pa1mKjjo/m4QtHdl3VarC8zB73us/d+YQt0YPU2uj+JfXJVd6vg8hRAHKQemMhNNn9dnT9gOS+
K+wVUolsDDsYXnPaH8U+Z4t9WZ2K/NJGfCg1h0okLyT+AvLi6/FkuGih4NwlQBec6XHgNSbb6li7
uIhtYPgTntIvLO9FB9YwiKCzE2QXLNdweX39m2P4xb4tx1hSTow+swgy31qZRZ3B/1mewdhbUtuD
jIZ+hPUoehKVOxnA0Eqq32s+q6JliAStuhCaMNc2/gZ7ymFnZmDiburQv/5gIniluDl6tja0AqAd
I8MI8JOCf9LAHJvPU4IwvJne/pRsWdDkkt9Hs7JbQU3KZ4e1UUZfhcVJW5Fh4bywWYi20DQppL5y
o6+YubXpZji8KAzAcFHCAditHaqHHapgctl6iNNrFoyKt5nRAeojUae0djsB54zjZNQwwuKLbEgq
q42FPSLaZO6ef5NWzn+F8KitGuxN+OXEXCcqLyKKJHJoUSRq/vZypSDAuW8/jOACbrgVDyjS4722
OkWFIiBA1Ndst/ETJeBxrNut7Q6uVTSf7zVV86fS+IF3XLkkTsURd31mbvJaZUMEtglEOSRYnj2r
mQZJUfGmefOnrV7YMztrqvDYb4sgWxrlyiLKcw/3ixqUIfEL3SKNZoRcp+nqzHLbEiMmjLXfCNWD
xvhVbvHKdlTVCiErv9js9IU10fiGNw4bBK+CmQbrpjIVCC8uSyE+iB+eLXx5/AjVR97w3PtqVN0j
kP03mfC3lApMY2DatVAySnmOdcLzZ0vxml/IOojikh+F8aaw1/nC0Lx8EXlOpKGlpw8O8czHwluK
ycKgTL04YoGkv3CRuKsw8UuvyzzyI3bq/wlwLqAmdBAO+0w9fyzI4uxAD6t+2VqA1z1SwDy5pS6R
kQuxn22KFcigymaj6ShzJyzQKM+xAHFKe5kn26txPSo7/1f9jPThRoDBHLNC+ksJXn+WNWC/kOJT
bE1lrhtb0nppQDUH0PzDpSjdC00eAJUJOM7WmkQ6LhZ4J184uavyobCP92N2mfgyLA6cqe/ORD9s
DTViTFbCgC8QBi0bJYNcdMNbhtxKPTXX4zN2D7HXG9hSyT9TUEW5iYExHTQt59TljX4cJl3NO2RY
IEwkpcqjdGLVYz5UpR9+Tr/2o7bftyaBcIA20H6q0pWK/3HFELMfwJEIVyuVxJRSoZyseqlYlVQY
uS5SeJbTzxgHeT/7kceDO4TzbhLULWx9ujfSl5ety0HdaYLI+H38hoJprErunnwieBsdZjWJNd4k
nqKr9t3eZKvlRC6Ia4tV5DHdhSjiwzWskbyzC8hgyhgE1/uWNMhkQ5AnyhGAzjy6QkUL16Ymr9Gm
9alnB9xMWOe/emwbZhLfobi6c+dY8jepTibJMtA6cj/HKfWQR42v8OvVRk1vjVvYX0EFC1o1rpTx
YFSjzRUkvJb1Wj5A5GL7GjFvN3Hz0GfMzFAACZdZ+NBHhwo/ssznw/Ee/pl8o+CSv6VL91so0SSD
+lpGvXBHz520EfK4OUA20uc45PWsSB45C4SCtwuh2EGmXpX9V80zLHBWStsG0xGDQJ9PuWg12r7O
LVXzIsfBZozm1nuZKC+9aZRo6DXt6VE40FpwIW1UtfEOPRQ+QV74MZMCXxfUAPm65/gtUm6rQ7yN
Eq5mtKcoIcZT/cQeimcO2L7chjhNunS+TtdchFFbZZ2lW2xghiDWUvYePxos1ew3PGqcbMeMUj8i
Z2sY6NQXlv7kdb00lr+jazMc1nKj0skWm7+5RCFfJwvvEUcAYM1Nvcc5M1ZAOiS/SV80arTrq30h
xU7XN80STUpzdqtOvp5nI0MD+CctOSVw50TQ51kcE6IN5spQZKjyP2XxYyAhFO4/kuFGZ9txRPIY
VHaVrkOriQOPkfJyHggyLDL0IriegOF+q9a3+2WlvlVcLjZNYTwSVhq9R4Y+ri7lAAE+RobWssGK
1ah+bfhHWlVg40qqhx3JSaVwOqCwCEnWtGPnYBQIaw2NwhLH4J4gp8pphH/N0XgFVRJokmtu6O3r
fLmC6ZT60mjdt8gYYmZwD5NNj1E0nmn1KWyIhqgymKmwBn21gu7ltk1Ymxi6BiWIyJABZJY0vx50
CqeFOpEFRBiIjM0wG+SEBWu7s93g1LICIKZBmuIiZO0BtsDq0ZR4x5WwTcP1z3Xinc62btxBP3Wv
VkFnToCSKByWkZzJh/cZkiHl66YkafuDrNvAcjuXEq/+lFFdBWsShOyBz59O6gvcWMkhV1otCPyl
WfZ1vR5cYQ/dSXkGP1w0Yo+f3qjaCSJe4MR/bqtfcRDp0Tp92ag8wOvitRK7cDhh6KA7tfcglO+W
2hq1Y/DbJ05PE5Wx0AMHuoHk3iEWeJnPGRvd4t25m8Hsd/JCK2bvrofgYJIqHfcmw7NEbdMr5vfr
X5BS347G48o5wed9KL5FXJBkO4+NJYi5KwHUv1VFpaphT3yaqiYTIy8OKlwCYjGYfznzkGBtVe90
YfX79xsqaaBw6ZcqvC2W1xzPYVArAku7KdzjVoxN0bVAN0Vo+oNANQ8r7WCmKG9FhQX5hgexRYRc
xG7ilczmG5fe5du/RsrMokxm+rV8OWeYWq7XQg+c9dozOKL9P+xnFWipBC5kHnUw7TqU2easHhQR
qeXFvo/ux3oW4chV0Ys27WcLLwA7AhdAC4IP5iBx+gsZ9Yx0WyYApTz/1QaimYghC9jLZ7SJMPjM
Yqnah287/w5baTP+9gM7+ejqwZmGJH9eTCtdG4Phmp08evX1tNxIjpHChwWVQNDTymFNtAcyE2Xv
Lxkcd5sOGZgJ6TDruh/ukWmoU3CIxHwNv8r3UjJvOIeePyfOMPv1XUo7bJDNr9LFlgkiyb/BatHV
ea3yNaBhFRQ9tYX4NyRDmVzdaIF99EKALGXJc2LgtgyP5P+NXqyJtz6FVyHa3zC2Y+NWSqSxnDkP
6x51pQQkY4LqoCkhlmXAseldeikS63L21VkV4lruftoRxiUfeVQAWqFfSXK0flYz6SfbTAcIal76
yhGrFQ4079k1y6uHAsJRCv2grq6ntALAz8qzsq2D/QSs9CkKpIvKsXdCDRVua0pdl6uHDicaGaBI
stp4oZAvV3r8v/pSsaHmManFe460rBK8K17gw0bgDeD39AbxSU0GYIglRpIH5b0cPPCJcMv0i3TO
u6EJ/OxdLbGWj/IgN3e7C9DOqnU7pqEX1gh6QQmpOgS8ix0aHuLLLtMmDveH7h0VU9NWnLggsgkP
8YT8phYO3n62WnRE2dmwDnSi7mZQOQ/QcXrz/tepTsxrkyzfRh/TFrApsXrFLT4LTCd6asKm+UlI
Dv0Z+unZVFgpZ8oqvLKqkKkF9n2oRzsjSXTTkUXIYcmKhYu6EU+J7Hc/+9Pybl+J/F/xMW969uFN
HV1v0R9ByRo2Ooo+LTlNANpJEZf94leSvEASziyUOlhrjAY5zjPOO2uJAfoW+5+Avpz0Q2oyPk14
3ZJ2/s/LbQZHV0Pto+mYGi+jSHrspN82DAiPClYfW7UquMC26Xd40GljYmBSQ9sI3ptuQkHBaxJ8
Hpbs55IcRBDOyMZEi8A7hjYp6puv94c3xVFq8zL5OqCPvy2irFsnfjBVPivbDl9RFUeb6tDQdIw+
RBZxf+MDicsFF1CMfWtZUFzjyA+FJExxjZgDLRV2XPQJ6UxNfNwwxeono7vajJe7FVY5R31GopgD
m2Rg3a1xPjXim/0Sd4yWpNyEML+udSwA6zUEgzeLzaswf27cnCmKhxIhDKW45v0DjxfJVAFtKEPn
AItNaYG1KBm6PysVXKeqGMTAc6V+IrgTydrAtUKaq7rmvLnSSZH2stT/vRzkF5Et53QXHvlZEWct
R4RCj/Ir5PHFFyJeY5IFiUqTdwQWhJ3A2rmO5N+zftl9zLWLzY/DX3xvUOeOyCd/eExWfgZfi7X9
rMWbthhCJG2KtButw/l/pzkRJfeh0fa8QJfOlT9SEv8HF64LIUtAeKKMzh1vrVybvjm8V8k7Aq20
vhFXDwquFIMjQiWWyWqqM8a0iDzLqWUU5o2GmbZ1BjYIjdf513CgyWv/ge9aeqp9CUJbXaz9iCph
MP0qrT6pMSJoFo/pB+3GrLN0pmuifGW6Zydd433hGLqs26xHNQ/v2Fd2O4ZxWeJAW8eSknxx04s7
iL1sBb59R2pVJFwatWha4izpA6Gxa9cj/YazIgzlr5s904BKo0uT0yWsYhoTInTWCRai0LQNfhFY
dJPXB+ab3Z0JUHUlGWB3tGAfdWVeoggpXuEq7SJxEYmdJZYD3iqfvDNcD6IXTdU4watP2JUwGML9
yVc2D7+Ws4xQ7sBG7TjY6Cbv5WiVQvSHcZeYESf5Gev+Iywx+d5D9JN0nJHQnXSq4fvBD+P3Y6u/
epieWlbjMANP7TT7HCcA3ujzmFlT6Oko6t//WCuTrWT6s8hJYu7jOVeqKns2HWSr3O5eTuvJ+LGc
ZadaOn0NtIecnN6Y/x3lk/I2ZvyD6ruCkQkA5qqBVTPVwUzT4hcfgG5qShZxazDJ6N4UoRigIk/C
O3RvVIhvqTNrYyBBCPwOUbqaofP5Qmez11gOs9OjelJOfd7cozRDBC4QPka4ZtfdZB2tbO391Yzx
TJWZrP7U9vLV/lKgmwul3KPlvHwjSrL39hiTpi9M2E11RqMesFd4RKdR/JMTip668S8xYUMJuLPf
gFhgp2TLEI3N9c95lNuj4UdXoz4L6NKPppvJGF5TFzBcX6nZQK/5/1dOAD3g8d8giaC8y0xsUcys
8CClZ8AkANF4ll0FHw2UljEJk/9fHmVisr7PaT1xtPVWHNhgVwfMDsUoWDP6c8DGeWjI2ZX8LElj
cpxtC1I/0xtYS3Bipp1eee0BDsyKbqqB9jkHfvrnvyCKJNruJbfcUf/PLOe/kUng3pW8Hkb1M8YM
so90LQfiRgSM5tEZ0WsQFtFkXUajarjYWtZy0QTloqeDFPUSYksVzb1seYEZlo1mYww/2hfHC0t1
7WtFHRa+9Noq6XHv72nSTuOhBm605OIakSsatS+jtOk5Vv061UkfFn1po8qtNkSu30WeABB9wO4W
kC1T1LNTg8d87j+6B0wpIjkjeXtZi8LK0LxrD53crkysHigY/G9ilofzDhy01WWEDAIlV4Vb1WhJ
fx1/tzmFKIh3vlfU0osNMdFdU7RKFn2J9ByvoYpee/NMU1vPumAADQsCoblq+9Q0rLD8PA875/Xc
gT4vjdP+ha4cj6MR/VjlW9wxsyDXvx5gEZ+0stQ56XajbaYZ8brT79nhcTWqpbUicLfxNb5SHrDs
AfDv3HbCVat6OIKh9andCHpBjrlalS7/+XE2rUJP+z0l1CRCXAYLp4KFYdifqi1r8UN4/eDxbI6D
YngFdFV/t2XzO8CGhlin3yY6NlYsDAO/lfCc5F8My/1ArcF2kkrpp13cF6MMoqxvA0Oj4TN+XOL0
W5EILjeFr0+7sFlm+QslmHXs0gXxg/NUKRrdmu1cnCBoVh1G80mtDiB45fPcv9YNVk+R+uhp8+bB
TOQJVh4OrFfXc/DvE10C86q4euO7l2jXfklU2gk/a/3NZjxFBgXjD9f81ToM9BZrlZLrs5CgIoNV
f6pBl6sl9BlF8SeYn/c0dg3CMcIElwh2To2LEaFN/pAbIRehmtcycUtAw6f68qaZQZc+r05+wSbC
65Poc9bnJMPSA8OeL2aHAY7Td3G/KbI+rydTFGfAVLCB49vzg8k+2KkBt4XASz4nyHuZtJZCC2gF
4Fzn8Ag5zlzV7RHCsK0MVhA/HKVywuwfxlpizv1rHX+hnP3kkDZhyI8Pxd2p66XgNhsLbB34nFZQ
rD1eabeMiur5YrPAVtqRZ/ph4Zzz4SASTnMXZ7w7KXgNdrwA4vngqNzhzg7J5P/QcXWPAGZpcziF
AWhLarfSPWFlWg3QFbTOneevzkXxawsWSVaBphliLcLFC8K/8WyJbeNERV4M92ohANkxpo2+fa9u
YElvOjU3KLYRUWoQcAVOYLQ5CL6OG+1Gjh2cIUWKo/xQXLkiqSHx/9bOG6EF1qBOoaw8DvxxjxVu
hOmDONa70ncaInX8UOTdMvEoXSQP+fM71Lkr497AJVmSblnWC//MFtbBOUGBymtDOQOkUJIv4NiM
wHe0QG75SWXTC7k9+vRgIRbURpxtJSCHk3CXDViGhidLkzeR7e4j4+lZZ1rvfinTdpMuDfYDtK9Z
YiuuWQ3jHi1USgkRtE6Lp9SnymICmojzUVcsE+O9fEV5gngMik+Zq8F2ciw/QHQhm96WqdeSIOnA
wzMKsa6a1DhcGTAJUIYSewQnK+Ipu7HEnXpNGnfg6Cwvr7CqEYvAkZcDDjfSD6/8PkZni5omhH7I
cKBFB6u1t35nv99Mr0Ib2Iotm9EfCAarPvOT2t6O0CXBT7kwU02fLi46lS47Ir0APq/k85xQD679
ZLBM5H8x1v8Ib9kjv/mB7gk2QLBWTyl7pWslnJoeUFUsXJYcvzfGmpe5H4Jh71ZSZr/GlQONtMlu
p1a3wlNe2yn7+eKjTuE36xBOj0ERm5W/WsUuFWwM+RDE/ZPM74a9Bzg5l4yb2Q4Xs4PTnlLa03He
7FHce2YjdiYWfiqLQENzFp9qGZvCv2axB0F3wn6QjPv5ydC+zGYGyG1qfEYG7pUc3HM5zsS/usT0
L7chZnWKnK5Rk8gk5DuRI91QAuybTQSZt+dMSHZhmskusFYiT78YBTyt/1onqMjkM3vTEX8Yrm/w
zQ2qNLLU1zOzfPCGmBRk0lCLNP39tp+4MNuJ1O/w/M3EwM4AHKrYwXw1eTfg8x6k5VoET9UrutTA
ryBWlQlGmDEgT7PFoDm36vMEw2XZyYPLSVhcp9+rEgCt08KwbUfwweT6M8tPCjwFCxv9oI8uO7yM
PU7lxoCkqUXwuFijY0gJgQpHP0yMK0dm2FEi+Opcn3+Q4apUVsLvMvch9TbhY0pzrkp1oC/vtc73
yMZIuB6BUDkLuV9gMhxv2x8VkGQK/+9u9vsRGIZHOSbi5PYViXo8G5L+kWyhnlfnY+tqPZrDGYme
93YKteF9jPff6T3skHXopfqNXw6taUhklmIqg01CB7UkGWb0fEsJ7YbWdnC4DQojwyv2AjMPpT/o
vDQ80HnAP6UHbH1oy9i76y4krIqiSuFqlvPRWQXTBNdLKqZdRsAutrT8/5G6tRFTaLNNv5jqBhVo
SZwSUgwlnJeTn3vbs5gxUBgWxSq2/Q1e560t+B4tpK6ypsM6eExAKuNbVUKygc70GdRvbWKre0xn
3RropN/lX4tBxwkupp7ys5BLVdSeiE7pGkcC6V5ZH4gpWG/J8WfbGRXjzBtwYyY+f2Ysunc5Vxh/
UvyJ9hVZ3q1nolKj9QUdwpec37oV1zj4UtpXs2RVn+Ahgu/XQulIaNE6OYqCFueDqnFvclUK2L5F
gsOvOFfQXh3gpBWnuxakhqRbAYiE5LI7UMymdmvkwNvQchKkjt6F8cov22s1WFh+qK/GOGLrTOsD
BcaTfJh1RM9oxYaiSrX8/jo9aYda0sEcW1EFAFNM9AjbEJebCqwwfYr0wn7f+g6GGphlzvfvMNSm
WG5ZqDoJSp03iVrhD3w1v7riw3hEbqSWzJm9O5k6NZAct2klmGCVzSiJ1vuLjGOwqUqLruCUceYX
HAOIiISU6n3EVQP5wdGfzNfmR5cqZwNx/P5SgcOb/zbtRcbSdaAuJLlatBPGX/vJCURN0MK58k9b
6a13xa2R+a+WnT0rhmhkcc01UI1pDv0KM53HebQWs41pstfvdZTa8gS9GlEvUmMxQuYv/bmPjSvb
51F0dqKlmJaQXDv+91aR+q+yED5NNZ+/bkEMhHPR0Wg8MlFHvX7t101cbLchShgRSfu5mxLt0rP7
dzalSzKJ3q8FrgI6URB+QgydMdnMRkISrd/l3+DCDe0d1KTtXET5iKWXZkdmz9HLB4XfieZ/q1Tt
gmWebyQWX+Rto5IggYKyOb4q27GJ7uXq9wITMVNqvdw3pa/C1rYhGw4oAdBMExMQF3Zwp2aBFaFS
yolxIWdpYns5fWv+1vgecmBtva3eAfVeg6SiJXRnzuevM950wylndBw5qDXRM0f7U8XglNQhozJx
qJG2YFQccyPUPclh9GXv7LV+VcN99yNPuJbJAHn0dOqp0xca6kvCIdRhv/0zcRlrjxvYVVwDJQCJ
8FFXvxh1LcFFmp5+0AETNwRY+fRZjF8C4eGJQFcd1lh4pOIN8qd8k6MZKModg7JdEVFSNp3B7lpT
cM6nZhhc4nFTCBqzZeDfi8j172JlQV5YW4KMnKE2X9/Q8fjOKanGkXZhbmSGrgiK3ZvZJalQTSas
Hu6iwDow+nPmXX5nXxsXn5+A7tnWHx+pbXCKK7W0YdhSdWaXdatBboPhziwuA+KLN6w/y8GdC3b/
bj/4yWV3kIPOh74PjCHxNAycvg12xREs3g896ux+YXjpM2Gkgjbeug18IHnKbCTlQPQI9gl+cx3m
rqekjQMQUHgtwKh+gZ3nbd8KAdP2Y//6TpI58CK9vhopNvqsyQgDIbAsoCWA63MmUoGzAPfqQ/zP
OEkSWZWFwFEiRnclMx65iXsZWNRXo93USUIpqzBbNGLgyliXAgwSeJWV5lh7MOKfkhkL/MttgjXo
zm7JtBhraee/qxQ+3oMMQRGVKJq1Nu01LyzVTAdWhXyA5fzVWRCOjTt2m4Cp3mwWfxXugYU8Ll+6
d9Z6JPcKw1bzv+hmP8XOP0dZ/cVqo4Xw5cy2dFYagNdC0xB/0Edo+EUIwUccArrI3EgEk7gIUmJz
QRR/XAjcr9yBzJHpJ6L4vR9E0h82fVJVNIFccQ2w9KMegR8iq2y3551U/86nBnnCArFDBBLg5mpX
MD4cyLdRsYD5tFM5YD2pOyERayn1+dhrkXwxIH6Z25oiA4kZbRSYn0vxOgzjw13TTERVitQF9rW1
kWB4Z9ZIAfklPZRpSFH4Tzhc7zUGCujgvmErDunAiEXX82nJHy/nA8LWoLUpHyUpD2696wlwWkty
SyYXLngNKFQ3Aio5+mtsWTB/A8VZd6iJFSJ/2A1+6mF4ddvqKzEG7Zas6hUDwvWB7P4aY1AXdpQw
dotFbyKP4kF5vR6G3/vbzJ6Y4xCtXDmjvWYzDdhrcGentY6gZnmBPPB/9XzE23Zzrnwq9wPoECtu
qUd17jQOaNGotvYXmZFjiCcdixaztobtgHeRxWiXldBFKDvMa926Ds3FpxwICLSLK5qgBBRz1FzU
kGY/hE/erkdQZEWMIHa9dHfEobn3HTsTLY0s5Jt+VivV3pszCoYFle5wtwUJhiWY0rkSai+5qo0T
kouo7jmg22NvR9/xgKg+dIKqCOz5VutUnDAgFUfAc8/SUcLeCZpOX5RVCFS5ktFEOFbinhqjMu7o
Oo+PpHEgpDN2vm4Xk4cZYgOfWiLutvi1isnfLFlm7f0lYfMDIqL5Gn9ROqKPtUXqDi5Dct716NXB
Y69t9TrDWlZ4XH2Q+H/DQ1uHcIAZBnCZH6zSQl9SoY5Nem95GTrUwvngVU04/nyHTZobeCkoN0HY
dRYFJkaXuJomcM3VZi+TvarPMfOg6sJrkvwvf429BgStR/SP5cqUWOei2VWXnLsbPsm3l4NgsldU
C9Oy4uaL/cTaw4/D64NvZ9uAs5rr8QTnncrhtHT6xiRQjOLPAv7yzbPBVvIVVXELnWu0+kVB2qn1
/VN2GjAhV3KGKtgKICgImtnRToc/kTTq2HV63YNQ8RDSkOQkHrRdJtfQdOeDi+GA8f13kc1v8/47
1iRg56R9D4dtpUbYgkbjH8DauKM/xlCHC/eGUCdEf6s1aqD6oF+vfyH0n6BsmfmL6buuPshpsqmF
1l76Fq8rbhdrXWtEUAEB2MtjEZteWWFZoh7b2897ZlejSuqscwCo6E/LD5HkhpHXahuvI+yVioaq
FyBeKTHYZSjnXmQFuWs4DUSulgTrTddPMqhLTKkqIXn8HpJhOfiu9rLE44e7N6Vnf2heyPECfxz9
wWQK+WtCFW21Su6ajUkEGGTSnaJoow3oxpXqJo38M8dCrb0cvTJ38JfE8M61rLA4gy29sHQU5pLM
ivxlAUxIc2Zlj0ChpQeQRbJPV8TDcsPPzprC7MuyRoJE73SRmcKAVnAGjb0sds7UqLgny6FUJUdq
VLqfTT8m5ef38jBbJ8s9oVtiNbuE/RWrbWpwYBq48kXsLH0TGiUOwxpt8kUjtGQtgGpg7ifyjoh8
RUijBhtuFq72V3lzIDmDEqjNeA3hZmDXxC/ciRizmsSq290UJi/gFKpPbyCJm7rLTvyBJJrUXi3B
nHTkzeKgNzgn8fboJ82tJ4U+XLVabx+NsppsqYlw65dHZqzaRnsQ8c1Dg4mzonOHl3Ud+CnhUmBV
Pl/rhKFEZWxd6dxfirufXFLHOk6e72x3YgfyFsFd6XHYxjxXBCmIKCaWwpYpFVuT+kiIyPiTu9LO
Ce7bvN347pSVYk2gnlZGV9i+oKQ6t2hfvmOrywXeEKd6S32jq50GTLGdz6DToF2TEE854XB5RN/9
xl2wbl8PS3cTbmMKNZVys8PvVmDfnWbWX/iXvNoVFtto5hvwC6WFhVzPRsFllE8i3gN10to3goA6
ffg89mDaP+ZRQMfd5gLheCu8ZOnJIzdD0dnT4CprN5Xi8VF1+nd4FNkQmxLJgk6nkThoun5qhU+V
wXEFFImrKLQ87u8F83OdnkIWlTImpkvF4/Xq3hPgN5GroawrrxNRi5h9JfJ6fHR0lcMnJTHGPbCC
UQO466pFM7asyCL2KkUmNB8dyhvHT/yXojKuAgUD16CbBUOPn0HuFq5O8hByFiX7zIQ/X9xxQ7XM
sIullkaEkfUoWD+Kn8CMtoOKvYXT0lzUWOwhu2xFHDdalLmxv3Era9zjrdVSBwyL8wTSyc9jgbf7
igwyYrYWZRd8+8haGSy7H0HykrEl7MelDAsxHn1B9rCl1GcXtDZJkJ64tdzkYccZ0pO6ySJVF2S3
KopofqUa+4/UPeUUtoOXvgg+ygm1H9//CJP+FRZKqI8sD0jXFznFYprPsoobojF9sbXchukj3K5Y
XEpng9f9/t3rQSyaqq4vRbeyIYb33BcTTajYJEOJ8vicfNxEFvbvkF2TuzRZYOLugVifz2W6vEKR
MhU7pd3msjObPf6Lb2sCWi4l1qvuPC9skdhJDgG49srBSSxuOvJTS5AjNuepNk/1lgZaR95wZKKi
EnHhSVqGoi1gZmN8XZMNCzw12op85Ge9i6fck1pfS5rYixhMeI2hu+qQAM85uadOc+kNyf1DQl7h
q6hasD2m2e/JOEVHS+H5kiLeAlB1kJ0R5xOC7y67tYIzEwfzxmYrnqUKWpwA0K+EDQ0rImRtcqVP
UpRFRSttGMCjp5BY7lP5Zl3LEasR+E+dADwzMlMijjaN4kZhcMXGNRbqnTeEq3bRDz3N3btktsCL
/NVlPR0dRZrt+EKpPtVWyWc17fOntT906LqlMilmvSdnAL8wRkuVNmsLkHMJ4/FQCe+PcSqS3N+j
KYzhUdtki9b7o1zX7tzmC4iWGLcCfDPy6/QDdpJqcVhoY1935wqaLLQdKLRJBEmBHDAXd4xL+uaB
JQPEh4sUZaXroESxk/h0xJl+WikNsRQAMKshZkdgwXVu+KDwbMa2IVFrftRcFE8NQCROrysm0nUD
SZG8pzRyQ+hGtqVG5gGy+mG/YRoQnx4gXIqN4RnoNsV3FPsTtGdaZzOgGsJ2qxS9zU2eznlddnMU
0PSPgzgIGKJ5FtyhT736E0gLKwIWBtFDmLyggQsjFyB0Z/cHsltOZBywmQgD9FY0IPCp+5oI4TR3
ivtGQAZTdqrwAMzwHW2yGEkYAWyq3BfKJKuD0HkFFpw4RRoyQ3nrPxFSMK1PbKjJvVTZzNAm0wEs
oClLgQEUSp0Vk6x+3DmDkyCAUYAFZkhehP225iHWfz/L+4y/rbJ7BZeZ+LFdbcKKhqwvfLpWk5Li
CqN2OOdJeGby7Bl3V9ObijJwTX823M8z2l05u4MEfbEagAKt1RwHDNmYgPSAwC2QGq+6qbfWYb0l
BLvw964hNxOtCGKsOG7goM+SiAhYEU6ZdkezoS8cOHbieL9CNNdFvREkkhugeYqmRmXP6AK4iSzZ
nZeGi7sAOd1GXw7E8TShJNEff8RqDxCHn01m+A0yJtfn/TCTdTBFO38EPWSJq9wxiAPPu13QKVFo
mpU6Cqt3PNDRS3+/jsOB3EYFkJ7d4AUSo2kGiFv9YG0Y6YYQQ4dzZ+3gV2Zy35z9CVcorbl5Fnk/
4zFyr9pnTdaYVj423/OlkWtMAlgcGP5VXdhzswJRFwRW65aBKyo+RF/RgSXeI4ImzjF4haJ47u5w
69sm64qhY/D5o8JIbzoLkhovHoeB8NNYzCrmEw1zwli4idNja+btDDokhznkWufwJZObUKFsw8PH
Os5bj4IIAiG2noBo14fO1wS1IK6blIUHZHebaJsbgj+SovGd/WBXxQzmjJzjLH6HooE64LIU3T8m
nF1fBC4z3kyRWMc/I8qeIxQ5O/wXyeKu6vLTZgN9MOWta0NCTzye/NtiPjFLacbF6fi3u1iMNDJa
3UuJ7C2EP/v+9DFjn7dT8uy7ABqd32cNZVXWIj465VCVCUv/Xxlvy9AlqmAFE7uBkiMS/c2N5Afb
P6QE41/YyO7btStzaQ/zkgLgn5FV3InlKDnkPZszmDwS7Dzj3a7DSLqma4CAAZ+o+wZLwlxu/3Wn
E93BCEl2fM791i6yr8N3HTar+bUJkuFWegfNTS5YOTFe1F80QEmPkxxX4ue99EHLTR7f2s0U68FK
8ZyIDCSG1pXIjHEFjNUuD307qeFBpQ8JEjTpckji25rmFHXJSxIqf9nzbIu/pJk5Kcv97ovBXEbA
0VxW0ZZ4ME4muETxTRyY8QLiP5dJwRThzWvnhCVCXiFJ9CjZg225/lOuC8X6z/E1tXR1xpNSr2nf
fzzX1KCp5q+T908eglFzY5ig25T4xAQUEpRPMWQVM/TFu2Exmcq+exPWDqjaYcnA0yIaGjuxSutF
qd37g9+rO/KBbELetodW1KNxfAYKfVitkYw2p3/kwDh54GDZDWvQIb2n46arpfOIH4cjfNtGBPyF
ZMTVDbSjQdAnB6HhjNnQmmgxFGtTFewbvo/eOYOqFS358QZ8JDUeY3JJ7T6qnXYNjdZ7H6nLGRqy
4PF/Ohzq4hPrPXRhbYutUr8Bt1jm+WOOt0tNWfPJm2EJQV2qSHEcM+sYWBwnXQVFaT99gMlKF9aU
3lMudxvStC/TwHMmI6+GrNclodofA6NAqVx2cgeTlvt8iBYCKtOQolsMWtivfKL0k5FgcDFWrcpX
Ev3VfqLasJRAz5d8ywSLLztX9iWhEo1A9gcjDg+bhizhSzEw5scfOq/vcBU0KKv5BFbopobH6Rcl
FOqCRRZ2SGq2nzm4zz4tSgvAeiIjjaxuciqtp1uuXqVLf2/QCxVhdzLHBz1jIipuPZjcnbvY9Br9
U49X0TXExXKizkRGMb76xY78m+iIjnRBgYBuIP1AVB5OPComleTSMzH/GfQ71WlC2H46U2i5oSP1
20LrsCzqibz1IpVKdz5kpdALWJGEX14VrNdUlSjXJc9x3xN6QHu1hBvfnWg4HiLdtk0zH2iylON5
GccpYemPRvHjXBQTqfM0/A7z93eisyjAChzn5E1Peic0rFCDdtfLHRj6SfI3ZJQSjJu6N5q6rzkS
F6wQlg5umEezaQBCNqDSFBAJSp3He6l6boLeuQ4udHHa47iTXuTfDFLA8N2pgyU/Q/DHYdioeClS
IBvlydaUdJ9pekiw/qWkvrQgw30TStbYsFlelhvarhFApSdwY5uElYDje+xOf9E/KeTvI2fv2VLa
5bAK+cDsMsu0HlB2sf5+VzBRjMjJ2G5MhTbYWnNWXUGmIWmDd1ryj0NATSOmYp1MQEPs0hepH/xi
KzfVsLfmnRCMbPpBgPbyn8LiDWDNFpwAf/dKkVdvb7ry73xxp6GO65RY5jfMigJxl4NtIU0k7MSE
7rv/p+jF1xE0g5vyI6sRoA3N/vQH8sWVbCR9rorIJbmC3Ygj0Q9+WxBrmXBOt7CCkQKbHp8JapW5
XrW75dpWwqH561eztnTkh4vE8rPH0rFW1jNNArmblgccyPji8xb0jpUAvMc5Tk9d3W4Ktrl407/n
pKtVPPWK9QzzqwppYxLxQvu0MeEA9GpswB/AjBNXGRsQapLWlLL8nE3JF53Z7N9uicz5coEIbO5i
AnIB6mxIctwNU9e5Ks4tMDN+tMSaBOOC3lsOkhBvmvNjnOuS2ja3oVNAY0YoHQObjN2QS0PzyADq
nPWYlBRPjS3ivg7JwryeXsdT/fNfwMa65v6dClXpwNEphmrXdoxMavZ7w4yUtVDKDDOvDzackXy8
AHr8f7Xy1/w1zSwBNpuKhrj81Gg2qlgtnakpeZ4sbSKjk3eNIVEpUMJZHEfKIrSphyv1qyAzv7fZ
rcX18NgZS9LSnZfyWIF2yLYXYpch8YYdllGqc8J2p4JLhvPYRH8KUzKQQ774zDXwQtIQrY7YBP8z
lRoNisuFlHsRB2ifC8eD0VFKSyyU2z0cAS/YH/1c1O1oDx5DMq60G8evqA6SDjHzou8jAHmNTk81
nFltAhzFFG7j+7msJ2v/4qPYSzDDS2J61jLIoAGkKepDMRf5EM/mThyIFLbC2EIvxIdwLT9NbYtl
0FjYzbk5Rlhuk2Ix1d1jQzs8GhrpLcYUV9PycgKNZUKJWCaOdiJVMtRt7ax9WHmnABUaKx3Y+5lc
9iZ+6Wh1Wko1tyzdzJiPo+tslDmG0oYptzMMaMRouK+VYUzI+u1KWojY7uBfpEbO4Ed4PMgt9FBy
0YtYKah5qpdFGx4eHFyrfuRgP3yBacPv7+EN/wvrLwzgDkAm1Kssv4WU1LSUlGB2SeBH27Ya/Cuf
x06SsP5BmRO4kywEb3lonyu5LRSlO0+oEbiAd6JohubVcQHM3fdmaVRva4P+9N1ndIYGSmaeVUJf
JC6yZSeytbCtaL8MIkAgO6dvrivywwZ+6n+6wuRM478zSWV6+Re1muSrRNXvTDDxlyBFJNLLJDC+
EEWF0yqV62bnWHRd4gYoxY3yxBk1UIBp/UT5XnyX/sbMsuauxiYxxkDVrKDAVilCDGh59ytwsw3K
+2ClR7Wozr+G8wEse2YtvOBtUTd1McTPYNgHuLCKl10Hsg+oVqL0UwK3YP1VpM7Ow9PD/Nx6eB5M
8oNlfGQDhqodkE12KRD7aqKZlYcJt5CRqmLP13h71fSbEqcENLw59B7FAMPhENh5mQ4nrhb2fCmw
hMHAtOxCWXlWoTNzSU2rM/L01MG7u4F7eLpXeBE/r1PrSzf2helxl1YfjrASD/s8G6H8CB6KAKqg
pGcoDA+HxSx5TNdKL3ZaXk8o4R4sltrVyJ7Hg4ae2xY1ZK2LVPHS8zjUpYQPRMx2iLFtTrbznVfM
Bwt/35V+qgPsRL1QiuKaDe9dOhvNDUSLwD1IsNe/8ggYkFpDu8t+8roCOLx758xeehzgTuCvNz/y
Rpa6Z1anKkuu7UE9Gzq93/sQgZj75wau14tAHhoa0DledDQOCgZ6gBGjAueZN8qPdwNMdehUKJPH
kY3cVHPFZYj456eO0yMOw4NF/erUmjreMoFpbPIJON9b0nBDPNPcRvSbncpy+thYhKvuyH+iW/f3
GenuNi9gAQpioIHbChGQ8kahJukCl7+3+6w8rWBn2cFEVHq8RdrAzK+bJP6CKuumn+tmuyc79Ke7
qT48G0SMVh2xCfsha5vvPlDm14pQNkOuQQNyyv11VYeZMBNPWoLqiFqqbl75WRIMj0bwmktOIDep
jRYqpXy80GE8kk4e1NZ66woa2lhDMFnyfLtSJR9YVA8iAq9h3Qpo7Oj7Tfop1BZrFh33K6i4KF40
PM5ieJif6YMJ4Y2CG1DAMsuXq56Q9Pw5yps5ezNa61w/LqOJlzTKAb4QEppjBmkd+ikk7deBECcz
ee6f3bvRwJkhhSJWwLblsBHUlFbfrYVtuf0mmtLV2A+0B30fZmAmOPUkH/CN2r1KUD41NMUYhkSm
As4fHitaDkJIpjMHz88m2VuXCHjFzIS5Jj+WceShL41pgY+S9wC/EG5rvQJXmXm/05YHFDsBdPQr
JbshY+SUB4r1UGC8g8Yap+bZ6An9oDm0Qxua55bmfEQNfEHtuBN2+WqN25LBjkoqBr6iHr0JteKs
afOiTUz/8ULN0Qd3V7dz4W8HPT/szt9m97J0zS/ti61/ZnzJP0MlHQ3iFqLl/KMDUKBOb5kWdr0Y
lxB0NnwR+uFo+DHj1EYUOjdUilnWVVWG0VXErZB5lvoXA8Q8vytDMbRZimpgKSXGgPZzBbaxmz2T
RTg88CsoAk/etTrkq3E+BIjdPnGqDiDA+gPTxI+Jz2X/LEbjJEmOmsPuimteuEGlnWjGmZp3b2v5
E4nJ4rzf44OvEkuJM1aWKGM/bTUSRTTs2Udq5tcJ9SyI5hw9sbIpjVaIblq8DwOwdFS7yO0Z5UE9
J/d+Rh54vsFGsKPgC6RzvEpKWsvGDzzNdk42pkhsEOwIqQNSbPTlOeqPtKBxWk9eVjn7BTE82TzG
iNckaQ3yluHdQjDWJNA7bE6mgd2xtPDbguVWbAnxsX+kCIS4yFrWKr7T7vQnPuNlsm3NAI+hQbpP
aoN/F8od/3QN4LWhfjDkn5OcqJQfDXR9shl171Uuib3McYJnRCph6ezafpf/XoofwDliB9XyaoeC
Gl8MkvTw2VZj2ZcYaqj7E0KDglKXo5DrdKSjUaXRn9OItyeapM6MMecbn7F6w1FwzdjzBNOtdSrS
Mc0INTTpW6svTgCI9JqiLJEXcs5DJFaxkXUUPcSf7gHj7kVaNHD8YAdIyhLqo0cyRPIReUV/DPwa
J+9FStI2jx0nF0Niy9U46OCdMlqosqTopQqaea0raZOGAxC7x0QJxmlHmmxDVLgcI4oK1i6KoyNH
yINUPYaZOSpSqjHyin95N8r8XsUx0x0Xbmnk3PKeyRWovbWR+Qy0zgYIRgB2kxv6d1MaWJgRVUWE
Xpg/MSJmoNwBAJL52jpAmE13ybAOpwCKZNA9SGQj2CV2b9AqPFX7k5Lu9ZVWFHrT56nH021q6ceK
o4Jw6fUEONbrLBD5V5mvOXLJU56dyLsOkfMCsvnO9w1MAhjJ8xU+Nuwo/438REWHjDy7IBcag92v
bFByEYWGDiR4JcUR+opqAWvPNAGo3l68xtZHnphi7STg/QKgTv6z4wcNklWR6tqwno8vLQNXsAH4
+DyZOWxj0fFOXY+PeapobkDZSZG2cu1H/+LgaLVE7LaaMqgPZ/CzJWNH71MbhA+wFjDXOLRuvrG9
/RuIIjVlTA+hOesrhGLZ3YCjE9Y2O7RVlLSIcb7ht56xEgk187zzDEWl3wlJ3XIBxMRmSAKYNjxd
Qj5L7vPxFhFCEa2qA/3tPilw7na3QgSsuBqX62zOY8hpoDL0xggMTmXom/xErpvdytnteHMScF+x
ImIkKtOplnAhRoAHoS/CIiKGCY+xSf5sAVfmaBIyIInrCiGfT+VccCKHlFzugL5SYSWwyqleORar
1Xb1S3XyihUI5/CoQO0Ph1TgmlNdzL3guxfwoWJHe1kP8TheaHZVRXcvV39Dn4sxk32UqNbUAnUs
Z/Ts/l20MGNxfWCX3UfVHxvscF1yKcSvBCBaLK0o+KVTIgy4snksx5k3sz2bHVau49tUTeTmVP/0
2ai2jEhgDQjvDvWnDE2Oapqre8XYUaAh2joYMpQTdLlFonE1s7cmNP+fd1sLMYgBH2GDYoZP3sEp
WasYkvaJ37FVjuO6RPtDBEIA9G9oTpjoY5jot9mZwN5zCnoR3W8r9FVT8WA+XW1YD+wShaOHCgWj
zaZRvwhrPeTLOvT03WxlQcqFygDm8FEZsXYTYUzVLlPOmDqQqeza8uaRNTWctZ7n2twqNJaa9kpA
+51jM8mEevq/iVXBO0GEpo4yF9WlQMA+WHAnZ8uiORiCdLNEJi3IfE+EGJW2JhE3EydpXOspxNHP
Ht6tX7zyjP7VIbszyBoi/On6cgvmVeIzWQtWPalKrl8D8W0/uWuyv04HQrxdDewSlJs2FNGc5oRO
rquxa+u9V2ycoIKTKKuXy6sepYS5gKcaf0V6+g6tz8Y+TTmypXdemNN4jQr3SE3C/UVkyBJUDm2L
Q17rHZb9sUG3OLzHdZ/nqEVDHeXsAMR1iPToPIztax4T1h1IESy6gK/CZzJyF5RqZlDj7lLhM/l8
kE/8/g3Om0V2lWONmFWk8LdPBMptkBy95wgwLeNTV0VLmmgDtoLpSAMTawKPj7t0TVdUngoWhJRQ
E8BQ2bHoHYfFaHIEo4gUHQqNuWKYQAucMSOaYsr6OrIyptm8FBuEq8WLNrbidLt1ubdgdXXS8rvh
Pps2HhZMzEeG6SGN9j+1byYQ9f47ULCKwbzK2I67agUsR76nH20vLiiERjqgsmQt4NYoygw+sLm5
b+nDCiGi7FgRQuruF75CmG98GWr2VJt3zKQkrxB2VWvsl/E3+0P2UAevLvSUPHOzqZTp8mdW6OgR
75Olu6OcEWgrgHo0NCrzSMPMtdoZmnHBgz+BHukUK/oylqfDZwldudz09dc4PgjTWWXvQrCQKfat
sHBm00yMRSyiM5WjxzKvRtkRvB+FmAbU37pT0HA4Lz7ZEg8Qy06OP+n1nHlUeTqShRx0RZIYa/zB
EzrLTbnnLRdveN6UTJQU0bYdYiAOaXSeADprZBJF5fPDtE8Au7wrpn1GVMLQ5VQFkezXm7UqffZH
JP7s6+BENzAqZNhGVIXgue0pGPyXLis9z3eEHvyx9dBRu92T6S5/mNihzUwssiM0T05L7H5+IAxR
XsHpe3nuqNYyIFE6tReQo6gV79Wd/TzQV+LqhQgLvRC4H98EKjOa/R7LKAj0+4oxQdlGUwwrV/G4
1JSKy8BM8i0PKQNieLqaov7CWJrrI4Jv/h14blsaE+5XddzLe8D05fl8zA6eGNG55oAEP2Y/uSAG
4lGbMOBEKqFUGc2dUscCMTiUWhPm40xZxqhm6EVgEtxKG9lAMPyEU170C4XzkIV4BEkYA/2CYcne
WHJLzAdTBz6HIKPnn1BM4EQZLM4DLBGVD8FN3tx50s/YoISaXYFrtnKPMidPrFo7jEei/fkaM7aK
NSMlqNqkekLWZZzBKTCiTCHUn8kOS94kuoODGupfP97wRqfDgSmn+MLA9NzeS6MF/Xm1gcg0cTku
QnrxH7pOPELSEG88qyIdS49tYIc/QN1AsLhWQgjve7uyZ/pqiVFLqU8bczZqyEU6k7UqMHPwgX5B
/wBrDkVLFwe7r6lJCB96j+a/RXOKuQp8ycjClAVd0jS56sf2EPIlnqBfSoNSkgnsodIyeVFWSNYh
IuHC9qi+1Es4jkN57VHnfFleFGItVaWPYYsnBLyABCVpNnHeit16JKwEKoUj3KIRU6Sd/np/tjJY
LvyrvragvKsyI2vpA5V3o/eoTo+BLCclnbno5A0jwqyxAr+u9YtR3Fe0HnjoTwe6dtrYANnxNiJj
bOAXGdxQI8nVsJQuksgmzwuP3lkGtg8svC0CYj5b9cZXVwhyjuhHDl+nZWROh0UDt3HxC6mlRGAW
3aU+Yicdm9q1CD1HMzfE9X07tf+Yt2Herzww10/1AMc9U4jGa9bZG8O8H3VVpFBBvC1DY9J91eIo
G82XI8njOEbtmYFQgA9OTE4P2IlEogjYO6+KiqHwQKLwqhoMtMab57F86DfXUBAoFnzKOBOXRSrl
vTdtBNDMRebCUBN2xHPzQNvOaOR+Zn8i+ALEGejPTJKy2Cwp9f7PydydGHIhyD5Tc/p5mepBe3NS
fPHZT/r4nnldtFa52C1PayIAHBZxSO+XsGt1YkU+SXr/FQ1JLT9KcNwcAOtIi3apVwni6gWx8X+y
QwZVrJo30kWVuMtYa/9Uu8zUVQj7090o979HXBShx04ZTex+QP+G3xZRx3ITMYIywvnAiibnCg3d
88yquoBvWD2n/spj1ZBLekfJyt2gfSl5LdBXIHEQGp9jpfz6ji5HbvbsSHm1CRcQUBcVDKPmeJmy
3LLbswIXi5Ufav2yvl8DU/4OzCP0WPW+o6rDQZjhuSb35m3W97V4rFZDx1U9dBk2lsHoNKr+uj4A
umhsqKI6ATmlBDjrODLFXKyJpnF9Dxn0C8r36cMT5wuCvwsJ44CCEgxlyzWUX//c+XXjzCzW/GAH
2YQGc7wDRXCQEeW8k8kGAWRqPhs33r5iHB7qPuVBx57NjNFPB2wq8sdrniiqniQ+QiANR5ZJYDHx
K1eWP0vlFZVDiJTO+6c6KcyoyXm7r5cajQZcVUgvqIAC1if8lXEix/Yx/LZoWRAhD1pShvFyd5Tg
Pig2mkKhYipRpPX1eF77eZXozpr+uNjlgjn0q70qaawiD8G/Ds4Ra1bFiXbrUV5o9SLk2GN2T/jV
sSzy+F6vrmYR8fI+uvPVPC0x9NZVgXmw06nngZQeIqWgEu/iTnupQk+Q/mjc37yBDFHgpIfutJOT
nEXOlVvkI48U8CYetqtiSn+Z6WKEI2rFrlE62RAVPO4CEvgPU9HYe/uHX2dvykG4aFtoI+4UeaqI
8ju6oK74IcFuH7sOh/UZGbmCA/SwQvyj49/IxNTikJygWDrnN0f4PfhqEkkpH/mJ63QfifjXlJMw
cHaaq/YiT/gHgStEE+tV7afyWDBZLYwiJuE0hZWJYjOroWctedv8BSDRG9mMMAi/EzgoSfS07nqH
53rOBQQiWYOdUdADh+jetKk+/b1qk43RdWmmbZon8fRSuhRc6a91Hbjo1gnkrYq6ONs3eizlGxqZ
CvFuLCYNP/stzkEk2o8xxOht4BZwdWf55tTNDl2t2PhfhoilWJbJv1W0ifkYppqgvpzTJVbGfc1d
B//6BSz3c0szXwd9RVxAE0XP77jCwt6DCnveqyazgBDrsblxeUZ/CoK/dMxyAVsReWHlDDjsJ0fI
4qANDRBg8oX7C61TuxsX6H5nwCnMBe9LRtL2U7KZj1GnNVijcG8xzs//dBJid+z6BA4dk9QrnH/E
iIWrCi4D+0ZWcTmdPE8+7sCnAPMEp/EGzUmeK1SF7G7YMP2iZAD0RezURN+AydOgJb+wVMw4LoX/
zbzHztoDvc8cPx8aqnZPKEWWmPxgyXsPdDgiRPpxMtodG5F09BcJLb7uxnd2aaPK5TTi8dpffvNV
a5IqC7wDLRP8j1woNa/ADWRNjEya0T2Brv+UpvcdRgrbdVHlAdh5VxjWfchUj/3sanSrKSXZxMYJ
51epovq2+Gh7ITng+Mj364X6up08UJwkAnv+vDfxceSnmKBlHmK0BXbzrj6vqer1qjsBW1overkX
gaAhWG8Vh8lNpX3NsLNv1SToAVBg2/X4s93TJWAyNEACvYTojfGl+AX2eDbHrVTVd6dz8D+oTytQ
jGZqS808NyeonPW2LbQGHMMhMQVZ+S+bO9YEESX4xCxdJGQbQooSpxdAv44tKgdNoIGPW6C4zggT
JWF5hZr0zDLoanud3SFdaIRhbERc15hpFU2cpbV84Wz6ZO7cJJy4RnwwFXs379AcXZ21TZClZFuE
hIKMKi3xnRsb0m3uHTtIhThPLW5MGgB9pOlpm4wuyVra66cE+ZFXftAj4jkwdyEyuOwzAQHHerrD
6YUQy/xkwLR1t8JgqRK3U1Ma5rBVhQSiyviy4Ru/ii+FRmeCtpqBifGnyzFWG387QNf3otP1ZHL6
QaP688tI5CuUct+rdfFvqlpAGqrlxb6wt54TnBWQN22YvCe9YFOm96n4g5b4RZKSuAvGF30lh0DE
wsCDNcVEp5mUgEadD8+tc5JEBgVjrMpq2Vlokpbrq2GJHlLqdlaUbvAr8lQUiRLepIO9g0LY6/n5
Hwc/usEZebxPSwyycQ+oweVphQW0K2ezPGoh2Q84hcKoe7J05+f7wJXwoMxx4d/OHh+sRI5Gp1lb
8R3TDCYaTldAN5dlIxw09G/qCfIlwWA/ONK51vtrAVw60iW2Vt8BqQLt8fFosmCbB7IjVhpdVRJ8
pQnNE5ecK4NtkprSjzlrdAXCiOa0xcKNFCg63hEB1Bzb4yl2N3mqtuHNB3XqAnp1EvA1Onq69MoU
JGF7k028+E3O3hb61deMIOsedWA+7usMNEDCWzgk84V/fJNeOK2S1MDdOLVSNSCCpmYtyxazwe7t
5nVhqcfzKLFW1xOw2yJWLDFEXwl/9gVX9pZzAHmyHP7fqW7iYpomgCfXBwkqiz768Z7NajcE7hpR
ElUyzpkwo0xKjTpE6yY4Zzk5DfLUX4uGQodqVx2o52i6I6sWpGTj67iTfc3YT20iNTp1ymUbq+90
ufHKIgS2oBAflsukdqrxamjgQGmta/wZbeOFjjEe+O3G+bjcRCUxpqGih0ZH250KQZV1UaEGwf3T
k7le9rnfiLvY9X16Bhfy+YLCFYRm//tHII8MxLKhYUXgYplCRIQPSp6UUfj9AXJwyVGDOCYkgv08
Dfha0Y+Jwml5saZcrfdGFn575nB06Yy2iEeTe1E3LrRApD9k6ltyYAA5iHSkdn9Yhd4JSxd4S1KP
SrW6Pzq5dIExQGR3qVFKijaWDrwmiLTiDQqei5hD4wWrr+5nNip/SwtpVak+EHBozkXE4SO84DUO
D3NB0uGk8Sra6zrp1uh552++G171OwKaEhc0eBjn0bGPxVUV/cyGgWNqdSoMemn0ot9mr3tgBIZZ
bkmhk9gfY6WG5AdgBlD7i9i8C7qRCEgBegriKUZaja+U+rEF/5V2KioaJV+ZDxaTozhUDtqBD+up
mVkHE71K4Dhf4dlLzsXSbPLfCAT2Mwu/qYGRXWomO0x0MHmas0Jv6YcJExrCzwjjDC78gEh5KO+n
9soGuRhDgAwZT8JPwbZ/KRudCA1ninCno3f+Auws0rDzORMCeEKznTvHX5ZACQb4Xd6RID8u7T1Y
pFjJsXOs5D1BvnmnULSVjc/eyW3L+/CLlvTqyw7kJ3GRQ0ZtmikRfRgCbX1Y0Y4RYcGA7g8RL182
xh337Hy1Qukw1Ic2n8CJEAwdsYHy1PzpGhxnkC6JytSIIaj7Pf9y2bub6V+FvCihsAWVugC9EWL5
Y+vJ5D+waakHbyu66ptzvdsLi3L/XriRVN3FCnj0k2EVFamoEf+0XBuqiWzb4q929q9Qc2Srn/g+
9vOay8LrjChCCuXtifltVSC6OuMf8pvFe7dz5gweFaHT9/SL/B2POsLXVtD+Di4DCnVXuMW0c5KJ
zcHipefW4j6H9q0p4RNoDY/hJjNjres7JV/5AKCwo9hfV5Srt9yI4v/u5enV8dIvM0/LvW/h/5iz
Lq65dOmB3wiSpFFNyXFQwWIn4VfiJY4x+8cqyhwT9s9zAousj+RGT75yludqWME0fbgNeocysxE0
keOjIHUBJVRLiR8QEkqmS95Tz+4l1LyebrJiJKAkf84GvI/QBaJA+9SD6wCWp1oQc89O1itr0i/x
MMaismddGr5etlxYrm1uLBzUzuNinVKVkraSZG9jfc/SQ4lZf22h1itx5jjxpDkBC9Bx3y9qPCpJ
AgRUb4WMQRhTMF6HItJBbl19ia/dA/O9ilEgPWqQssxIk22wS99ZWQejZdAJ5JYs8WnZ4JbbSw2V
A9fcoYwty289/elO7JaLIZgY+DIi7THRzspxI42bggVyU3JqubTZDAH7aMQT5SdsJGhGqu5grv0y
BrVpNqxJSQ5gOQq1QisMnXi78gQ9/QVJrhRsEB2aESqhLQm3HBTQsqb5SCKLQ5AjFx6/ep0wsxeC
uYkfkwQE8mnLXmCro0K6V9P5JOGRxyvt1unX5Dv4ey8JKZ+Kff3OXkl75h/mfh8YXys9fJ/vAqH5
n9RMEhczA83COK7Wwk6AMJUZ4mKIUODJdOcu2rLy0AWuMRVKO6xKu0H/+NkLWKesM5oU7RLBdocr
dmTzfticf6gBEhw22EKYv8wjPFsvU5t2khNaaaExMntEwg8Iu0eTmpmKeI5BKXzetoGSsefEc5D+
Klv8CN+od1MDQwFil3bFyjN2ijufZ7zlVFrlsSaHSJCVBz1OLRn6qSTZpQReYN5dKPYQSJoCOZBC
9mDOODIf7YXI8mq/nywUPNy4MsD53Lcqri8Rslm6ucd7p2BjAspf9n2TWSpDF5KGG1cOuvWoiyoz
qkGgX7BnGN1/us3skIFJctNSzgnjYmxDTmNQpbqXDXRgpBiuEaEy+EnF+eQeKtptEY3S52FhnyZh
80GRR0imUenXg7bZCh8iqBvvfp4ggTt7OFIlAoW5B4SUwmUXpAXaMOWUNG3ZLJJQrbfDsRCAehFm
hqn4itn3bVn5Lzgdrp/0Cwn9Il05snKL/V9khsk+bPuRFnBodxhFqsF4I8uADrKyDJLJ/KWAo3oN
EFiMCzgR2p6bEdczF+IOEFLOoNkKk4sYpLFtufpl8xWSvn84gVMifm2g50Z4HkRXY+HJvXN8iDnV
CFhOoyFECyI+/D4b4QT9mgpxyTfYAHk+cZMm6LllBMgUpimPOxtjCJ87hqgeoI/q9ovY105ahxIc
nsi8aNtRMxE4atMI0896g4UnVWrc+lH+j+Emj442oU2nm07rEGrJ9XENMmbEVNZLxTL+h5ErbGuk
yqEwWrgDfSsgV0WceI6couYevb2FgBxaoixqFuwPcYzJ4n6zhTOphD6KhrucVzEWp+v7pNN8Ghsc
tOWk99JZ3kVo65UnbFaYOBZUUmyG4le4TS7K78312gshDyxG5SumAintN2QYj0P9PSTmZLpehaxY
4fbqs+daRNpIP6exZCjQOiCltlTqjFj5Atbad+2BcYRMYW621PalxrQKjf1FVuYCMpLwW6dDGqcR
fRokbSpkneqEaGrAcNXI+CZ5LTnvSlVlli8M/1gN1IGk2XaTWgVjnVrEYx0sheVUIYBOArDifjQT
RU9lWB5d0VJPq93NBhvueNJj8OcVyFdlfqI677tfqTjkDY+rA5vIG/VQw4xfJsyxYoCN6U9Z8rYm
NLROiWpap59GoiBFVpsNu+/fuX+TDNQPXg638tzhhvkOJ2y0W+PzLiaDjNAZvZqqC6gpUTkakXeH
ROWXOrqMOr3yx5IKyJayBE+j9q8O35Q0LxajkEdvCG0AqkAmTx6jPBCF3igstbObiSlpnKO87vda
Z1858h2oipqXL4kwOIiY5UZ6jvGGTKDZdgk0q5VVURiQAZ1Ejjc9NT26c1HpYZ+NrYTHa45wNN/A
y0hKVMvk0doU4OWxatGoiQBD+BjraR+mZbZWAq9Gkn047KL+mesx/tzhIX9xJoc2xTKTB02cZ9w+
3vGo3aktSug1sE0ayPKeAMNg4H5Q3QmaYpoALUNUjnELwyQNGc9rFw8UgBom9grFHrtXRMGoePQh
XLKGD4iM8KvKSvTE1Y6I4nCBrouQdjQROjDvxaaqgGiAtRN9QI7Mz/qSiqLV88sSS6tIiU8Wbfso
atVeS1nL4pVss3u5ZcdIN6S0/Rzceim7D9baXTYYI927HERNR5GlUjOKro5cYCnJ5hWKrJ4WuJHO
CICsasTM/APr0BaBhHsU0Xnx8/VvV8mSTxhdW0OBjE5tHzt8blyQE6X9WsenOwjvs8fZXiL63II7
7BAj7r7CHP3m+U+1NE04j8CWRu/B7IRO7GA7gypHFK3n5zSWjFOniIA/2F/PC5u/f3FiYtqdJqlg
UFvbW7ItaHxhrlFPMwQAeos12Id5r5kFT/E4wFEcOHKS7wfgwXlTh1ei+sIfZlcoDih5AJsN97Qn
6zkMPGEvBHyVobjut9e2Pvve9StQkHSA8Chkb0Rbbm2IGJMVQCYByr5D75YFUpQa8bBUIzyDYwup
Gajv7BROJESPYPptfQNsxKYAhc8LNjVexmBhcNLbI3j9kCviU20V3na6L8AbsJ+XgsE6TtGIYIXl
q4LjfOXHa4E3ofZ6PffA2VFC4xGxF+jQETKxeJ6OkSz+y0io/b3dPimzUDQ3SfmJj+wxuxuCQaUu
DlFMwbReUX74Rmjkm3+9SONFTMG4vGoaIIqLZrMPQA+zdnjGF8BjyefIVcFh5Z1VvOIzGfQApwma
K5BB0DJyRaGbvcvJ8zWFLiFUbjKfMq7Smkm4iBRCJXtKJSdzQJJQkMhTCWeLfCLz4FqGRMsklXtQ
EXOY17TWqPn1e9w1ihGi0AXgBrFLNkUX9Jq3IsilsepJ4Z4kqwagLLV/fnlU9RV0dCDLJ8aJ+nVc
FBdDzGfQB5DYgLjBDBkUTt7k7x9805FSyehUHmNS5DfMAb92pdAncxfCoGdagH/rrAzrOpnRDaGQ
GU48/FDz8CvUXUyVwCj7BJIbMx47/a/4qeHFU+evT3/LtuKNNl1SjLgpLeXjOCDaQkLQ/NE8B8tX
y0V1spH5W55/5XyUFYei3eGWu8FGpzpjpjrc5wpwtK5BBJAKpC49w8ID38T1ZXeW0ZPWDMKZYFS+
Qn/3PIbrbynIwxLr4MiR05NDzDVQopBDTsVhpjr8jAFdmbUK4nPkoswzRfsrKbNUocI47R9Nqgw1
7hgG6d0RYUfHYDQYyCCaddTmXCpgBfUNqhvcl4YEoUbN95c2oOjkiEpP9SfHkZMEhPlOMpi+rdf/
qaxegLp9LrdorHlUKcZYqgVW/3b0mgQhBnGyPSGrOKCEj0XK7uA7zUOX89b9wseILFve0bvOo+hU
qc2rA8UyncTzLqHkHEOohmm4+OZW1ccYiio8PaafJeGT5n7FE1K4pnpGNNBpshPejevJxnaGVbun
wi9iFu0DiO9+C3iXaGTXPF17TbQwsvZiPYhkroMxrVza1CgU8MJCA28xoLKTmlMoK5ZT6uPEaN3V
TJuL8g9zXG0PJfn4+3kBF6msgn7RwXw/AeQjZToy7E5ezK85bt3BoCNKKUXM4PCRJrYLO2EEA5Mu
RY/EmaqzFtptDwuW+Z9EIhbOci8N3tk0RUJ3FoexzAzupmC5KIpNs9uPJ189qL19S9ujeGhTKCK8
BPri35qXpkzHZw+LkfQscHGITCjxOnTtHdhFXPy93N0P63OzR9WKBITyz5iLIvM6vpIXGp0RCfIt
5viYHXifS9RDSAvN8JmS49EdJ1jRCyaRMnI7J46hZwmkstyqizf7zvb1OTALX3i6OYlNKB3/xv7l
rYOrf4XLkm1UUp3zQdOcqJT6H3CXFEKAP2B7tNRBNTkSaWkuAAvAEcf/p18pqumzMJTxAr76QUgA
fxoeIbi3ySxhsbTkSZTxrFaKNdrAsSA+fbQ8r8aVK9uIMn5qDM77Uq5mt697cfoDaHFlv0DytaPZ
mEWJVYLZAj5LKtCK8dhNlXywLYcK69Ulsvmlja7wnifAFr94B8zRMNzO5Jpr8ZgkjK6/QBrlC1Ja
tpkQkn2THwcI9mRLmaLTee1kDwe1bcYMvKuv+6FNVz9wpQA0SBZ1U/U/B6mhHo9S2M2jH7J5XI61
CjCCerK2lshZ56hIen55S8cC8Bp1SVIvtXauje4+u7neiO+YvbmJbmuB6UpmxdArH5+lNdu4FSgh
rUPy1lPoWW17NOY6QT2WFQzYg5wgIBcdFN7P/9J+kVJ1xmitKomVbpanmrguw5ZabWWETBXOptAD
0ryXjQCLlqI2oPIrDi07s3/r1KVxnQeJdvDe2AD2Cv2xhLcvDUhYGSw6XZboVxlOZwv/R3eGH6nN
Jv25CWWJZqSFGd6mloFj85yawL8VPHV5syk4S2Goehz/q/M7RrOvgTqPaXfiBthVA+DiPH2X6+B3
872ClDdjE8D4tFllwDw5xdkB7Zgn9sKqBrmRvBt4HCLPa6+9yEXPo8NmE3pi0pi7Pnbs6uj1q1mm
hPWTBK+FjmonOFVgomYDgnAR8zyMUXKq6mahCiiASGLyA1vQ4fAi87b0uzshhlrZSZcNheufDroD
C3Yg3/2K7nKgaKoxGOi8sH/OCUA1cefqMG4KfwMNzeDywp/xgvXVZhfAmjG16cpHhCPOtZGoQeYn
Zxh4Y+9oDWmvBmOb62Ufhb57K0WXNvWqmKG8xdg/NCik0OblDK60/GfptMWgjWi9Q8jT9an9T3kD
vGK/GSu0FHwI4uD84JT+UtNXY4iApguyC0GB1wqFzniCY51CSS4ozC0Ztl16OPfBDMRRHyfMJGtY
p37EIO6RxW7vmqFCreKiY6MGQOOs2Q4sIYbaOLOOiBalDlPiv1OS3JaLorNutaAcbpIwDjfYmKQP
Tzjvynjik5vNLRvg4+2r48c3nAolSzV3OzNCegaZtNDA29fBEB8GXyXUnrgjvqsF/nsVhc36YZRh
WmwHqNSMdAZxegjxowqZX3fJUzxBdKj3keJkA3515PFU7GxoxIsbIpvopj9APTPcqwQchwo8TPed
p+xUtmN/u82Wv4OO3ZgIGdAtftmt6PBxxz43dOFixd7a9476BSlFe0JnTSCe8zwVZUY07eK2TT8c
EQf5jJHhFsXBp9LIEesieiJ9fcHqZt7g34EynPnaJ1ZA1N6RUhH84YpfAKJqnHNQgyqweZWaYSCP
iNWl/LxMfKil+1i+R8VkMYLNrCEuCUMcv6mbkRqA/WpWcLQHxUVm9X40fZYt3SbvQBGObBCXswzp
WP4XsZXpe4LkeK/yAgPISEeaG6mAZO7Z4IEuh6yP4LV4ZVJCtZbCYkX9wicY1D+g1oK0s349q7Rg
tFWtH7cF7jHeOFEDRm6m+QTPg/+PlVJegm02H7v/MD9EHAI2wqejK4zOtHaRkpgYAhcoXUsgIwIL
bkvBtkfsVajFw/VHO8sApjSEuR1NPda2POrcViKouZoRd4KAkps+7bB326e/YOOijnsojCjImVH/
5g8Nv7b8QPHR9yGC5WCMW4ZnCii9PfGOCnkdHNoiJdo/OUQwFjRwKw5vRdh5tePD6ds5bYuvAGH9
OlpRkJouUERdGhCE/b2sznSWf2vftiGT1fypfFBG2QcCVyhiTcdk+Ed6CuCzvfFeyecedoxtasm0
NgGhSPo1F0C9PcFyGcSg/yUmSasjAtwL5mwUoS1/bjK6BmcdNRjI9drZoFmhuf4Y7DFAJhX9SPLp
1PQNnFktUk8sUcUTPReUTdvrBces6FNziRAxUoZVfx0uLOIBtM2GBPkVbfn6BUjFA5FquwV5SBpU
8wVBO6ysiitNks3qd8lQ2GgdJzjQM7GmjB5sFh7ZOtfMMkEZPkbwdBorJ39JS3/2dx7G9t/NCAnK
lfwVF40fimogRnEmfTB+Lxk1fVmGqggKPYH8eS8PxCoMBL5wC+CJJ3Bnr0agqKE2S8GgOG0fsI48
gXYfCKi4DieGqRu6+msRT2+zJlfRb764gSQYjNYTqhjy+Dwot3+O21NgpFtcNXSqW6Gfd0MEgX+u
ecNQd6EIMcj/X/WHgY8o2edOOJzoMTjgqrOXXjhuzG/aH1ouCc3bBa5DSSOpJoUrj0yJytfwLtaG
H+I2otFhEdfrV3bhhKRiah3nkTL4FAsnmKhae0G1vO+1wdeD3boAQH4jqBo8jn2+d29EZbnSJZ+Z
M0GCJvKkLIBIHq3Duh3qmV9lRruX9Qpq+sbpNsjnaogPigSZEkxku9VI3Yi9ZxJkD4CVGNtV/a+y
ZRQEyjadj3acsDOGVsP7MbZnijLestcLNdK3tNRXG+uLkJlzpstBXazYZDz50T4lwxxPEfVJIe4D
lHVkorYMUGdqGVOwDt55UqwKVTB8pDKDok0KgCmh/8qulaaHIL3NXDO22KuihM1C/Z4I3WMbwuGK
UP3d6pF4BiqfPSsY7fVB6f1m+42MZZDRQyZ3Y/2QapybYMEtPUQBk/xWNoSdK2MiYo+odtRcp5bD
TUOf25LWk4dqnUTjV3WFq4MkSBB/jgBwv1+ZFCUNYMGRZgnd/AK7VQeDQQIcJlrHxry9KU9tqEfI
C87U9bgQr0VprfEJeg5T9KbQf6IHbvjaZHv3xdRZiEacIxV2JCq8gNwdpa7PfsziWm8biAGnzVlX
Oz40MUFejMcCYNbSReNW65qctiN4yjyAXePzAVstevbNVB20zESh+CieBVHgmYDdplBKX0tVD9Oq
d0Qer4dqxnptM/NfOy4bp5wgUeVPHhcm4urDPIb6sVy20azaOTRlSv2H9WwvMm9Lh8mlOc81zKa6
/01UbPAfO7spRzRzCgpRhGyk+KaxAB3TI9L3bOm8vzlMCTzTNCCd7t4sVypUq5LatkmNgAJ4Jv/U
3Ts3GlNuhiaAQPfzhkUQuS4IgaveaYV7bQ0dgkI3QLQaJyVdABExZmgQ/uGaizIpI8XrnWePoZkj
5ssSWlowkGmeh7s/sqNpr2u5+KBW8jSzjzFX6iIJ2VBiiuqt0HeVLFz0Qi9/vY0PYMKXihxm/6Jj
dylme9QXuFKAV5yLWSjH7t3GCR/No1VRStDicpkXMyztDpT7/dFWK20C4vw/yCsT0hJAfhQVUFyR
A7Au/tUsGdQZT1y4w29GgyNNrie3ahAhcbXIBfLzdnHx/suQARH3cvVZlHGw4oJ87JEx8mp3Ve8n
g1KFJQ6USIvY0uOHec5MLr+nGtrXhmjDJbQbUik5axKD2IKzmST2JF2Wy9XZ7IVMpVQXYfPM/sln
SxNIt6a1jhPSEaFrmp9ynfAhNfVUlOgUpC2L6HTXWW9e4VrWBC3DmHBKcnWjEQdqvDiFq6Doa2QX
xsllXfaOQokhDXpOth5r1pW4Hk4OQxuMCDr+lIXVH1hKSg4fIgD+F5wFdyVbhuGz9gk+145PScjj
Nu4uZ3MysqVHAzWYTVnLFDMAElXk/qrOkaKoMnCc2YLcW4nGEwmaXC5uxlDrn1g2XkJSLT0Bu2xX
iNerwHjIrEvVqM4sAWF/dgEFG4cv+6QZSw3PbVDC841fTb8goKDZnFRbFi8/YN0HjLHn2A9GSySA
jMLqyTZSFMp/wNfR1yHiEtz4ii2KurNdhTxcGFw6f7u+1oAX7mRw/UwdJdN+O3F+mCDA6LaNE27M
8gp3VWtHACPWmxX5DqIDjWhBDX9M1v+Z/6CnsTfFgXtSDOyatTl021hI1pJXe+xtmAq44qYXSwpn
ibUgzWGKq8fUrHtF3qFlXrqvmoZQm0RhOYRu1MyocAO8IQZNvUY7UF8KDCHhfYmJ+uZJg21y7dJu
zoNyWcRpG21nXAFf5fN3pJV+6UVRuZvffZPGFfl6uXUFnLMJqjNeTZX8ZuyHHZ1XgLe9GlcIjZSw
2q+LGOHyuQKSss6Xw6YvI9RZx3+vQ8MHcH844klSyYD/aWqk0KO8+tlJM7iuhZ/KlOcGAPPjgJyu
DA82Ev05Fua2z5ysbbeESaH9NkACjVXOf4DB4NYk6JySDNx4wUwjf26SK1qjTnAE328w74jRcwka
fQWfXcefwuDiguniZabjJb+9CYJEF2IblR3vKyj3iVMJ0KGrx4MeZcrQvTbg6JuhpSu7pYK1ksy7
mz06CtfdFvlvD0MFxHxFGZLww3hsjAx97MxrhGd2v//Cop5fbljTxHHNjUJslK9nERomjJctUlpU
dIcovKApe8cXtaJ5etOn5xX4wiqCWDox2c3oGPNGjwZb1hqV/c7AtSSSIels4oXO5cbsNdkROcmN
xtpAJFknjKl3a+KJi2uI0/dARCd7zFv8PIuh58ZiPyqkerc+qr9J9hRUttb5oD+8zucUGA6GLdkz
uFG8WxBgjecJo5O9Q+rfV9dtrCvIRFrRSBax3MuZlhIhPecNMe9ConkjgX+EryYV6pDkV3aOsUod
d6MSmnSOR8e2nYJPZgM/WSbncezVNpzQFpBEQ33gCbu2/ttJzHAZ19SNcc7zSqfV3f5iAJL8Ur5m
p24yEm+NZnigUbGeXw71JDj7KFTcbvVVOfx3dh3y9bGHm46biMDYk/I/NgPxlVA3PRIjMw7gxYSn
8dISWTSOgvgWzhSvHXPNmCCs0w5FNAulCHlWEjD9b2QsiOMrwksN8NTo6mfUG3QdpjdPERJEz7fx
ihSHTFN0wqvD7/dczG3KIXOf1Lw5biT2k1muZzBdEiaV0N9C92u5++aio1ps6x2gmL6AVemBfgvX
iZIKJp7yLulRMV5Fg/vyYxTAwCDvRIRjJyyN5oFPCeBxsRf7VctD/JhehwHgecQqgT/fuRgPhMgJ
jWXyuO43sO2mGHWabEUGwNhLaekmtRNGGGDXVp/0cGSAferayoTWX8+9wtlnf1BL/3UhjLRakKAz
c52Rr8+HKpB+VjDvG0s6FZFEqVgd/u0QIrUCMr6zjzxSlHEOkT7V8bZVW7HDaQDONwy+G5By2eHx
lJC27AhY7F+dtiq83aHPUbPZO+/ZqAU14HCf78SiLdQBta1xP65LqLbNJpQApApSdQKuqlVLboMP
+tFKaXy7TreTmQcV8v/JGOPpzFbC/Rv505uZYw8kIqfWgpQFjgA2Fd25PkifbWXRgJQ2CUVq+D2b
Gw2G1tr751yyitmjywLstJm42ra71e6TqaQBxpiRoqntcCYI05B+HM5ezdtKmWR/9HcvhA7fCLvu
yZaHGd4cAwJcEc58nnz0NeL1sRc6+OTVm3wBjjeGatnQ+2nF17sK0OBHAGWXIUCb8h+lxw2zBMwb
eTexexCy6v2yC3TdVf12/w6Y/1xWaSaihgVOJpgEQJZZQTDYgro3iV5WG6keqAfMZRC8Fu1HBTez
5i8EZe2bMPuMXmNlB+is5XgGfXwK/uW2G5mnfLx6U4OqSAKkHRiLPG0c80ZJDv6BikqkLL/YlvjA
6M+vX8wWsn2IW3jtfqWln9GL6rdUUsG55MZTHHqOpsHNdFgyS7982V5wgWeANF9xvynmqeq6ZyM+
jVBfPYURg/7p2xfmRR83ucBzDhYwCVGmUARJhkAZLH4ya34yA54szNmXlHy1sdP699D8VpZQ56LA
c0kkwnh4b8rkNaNYiAbt7T02jPSxnMG0HcAvviI/Uf8Bi73Zg9/PCRJsUruIKtTewRYCJsNUKGtZ
oj+aW+90s6hWOo0EKbjoOZ3Lmlx9nSaXC7x70z8Q7CXAgCjySJs7GbhkL/oIufziAfut7azceswf
fhOy1MXu/DD8cbQ5Wbs50p1sPA0Qhuwus375yzoTQRimHafDO0A+Tl2EgyUHpYNXBGSRC5Ky/jAe
Q8C+LD1toDYTK8HUC5KuIIypI0tBVgfDYMaE5/Dt04TxK8IFKBaTmXE6HBSctB5YQog8ryySTQUa
yhkneThx9KYSbvumiiUu8MwmYmb4dtqPu1eBGVIHBX/saxvsvtCdN1RCeojA2DRRasj0nGX0Vezf
blA+D3TOXCBqAqDZM+L8MVA7tyzexzHF9oiLVj4NQ+a1MpJ+dS/hMmaGADwHJGrUoG2ERea9S56A
GBCkhC9cRRityZyQu1I+FmzxeuG0lmZCgv45PNFV7+xKT2yFhdzDM/9GjB3z7rFVJNpsB3kVlEvq
bQ86FRmLtp2vN2lnOLifhUeUQgEaEzbC3hVpg8uzTpzTH3brB7yttpbrkdeHhGzZGT/bgV4qHUkQ
LzIdrL2FdN0Kw6c845B6A1Kby/fvU+I7STjfZb4R3kkwbyiRkp4XIjScth5U3vjmgcsXZf3w+spK
/e/XLFPniGAJGyJ640ZWKMSh7KoXRHPzBhiaD5UPnrM7tu/HF2yDCxxXPVAP+B08zVe1iOLcdxOn
zweFZRM4CMlwyJcwSBrOyfum4bwJJa02AB8wPO/SAoQM6lA7LisEthP5Rrqrsgsz8fQ8qQXwUhv5
iKnUQMDwgUkztkEwxtJ64ZNuShDYDJLshuEns5sTL/iwgldxDwput7qcxUa73xqMHiqT3WfMFKwl
wylpXdY7hDI+yhVoxVLDM8BrBt70r/BL1Yf7zfbFKK729zH0XyeRpc69kc1MIX2+klQfg6FJWdVV
h4dl5eAuhRUaTqeAY1obOtl5O+KRaAi/Wvwbs3anqAv5IDvPV6XUHi4Pi0UFPkCpQEbfB+86qQ/0
420587mezomukRshif7HhsS3W/DQSa/SQxE+5KU+0rLIT+8zw/QIDYkHsb/5gNaHZklbgtaxxUxB
HLa7l6R2teyzQ3ZpJLruNYKTFilDB4BRAwPpGCZ3ZvVSV/l8NO4soaZKDypW5iaJFK7P3AQkEk1B
WJLxuR9kSfVc3vyXGB4dRDfrahAJVsXoLKXiLtA92s8WHh6t02jhzrN1gnmFEgFL7nPWxsOCIyBS
p/UvnXMF+tjWF7A1bk6SMPQEpRmR3AYbeEXt41f4oYAoGOq8yNt3k++3lTaXGcASlN3GQPwiLg5o
b/82+jcwhi6r/DenC+lRT3dcdUQBFc6qpkKxvWx1VjlI/ToGtJ+hJAtMnlDCoWp2RerpqLTBpf3n
ZlVDXN8LcM7fuBw1gPJnSLPq7sN3GsPtWepOds6bT00RLA/H+6iko9Y781ZtM7mkiMFbsFLdfxo0
oRXzqL0/QBUuqzLK/53cD8zRdj2eS+SNvH8tJ7re3EMlEWZLyR6N/fgs7rFKHRCwSPfV5jaUmaGy
B/BC0jkDj3IRu7KUuQtbxcpP1tnfxZyf/PunERZ4CzOi+iHJU1M+qwYQfansZc/NBrFeArLotGM/
WWhuECOLi4uC+3U0jxL5VJc42RI2g+8SzLoDKmgP7XiTwRW4Jl/hF7+FrdO41VI1FN/MH+sep4il
/U9ULNRrmbfwUc65MQXUv/NQ9v9ieWVjjqaeSHuREluIoqwG3H85HjkDQqaJSt8XqRVeQLyz/9MB
kwibQ9y/2NRDPT7VPeHWIEt7rBWsB4qIZE1LX+iSAYF/cdw2EvlK17PvnxuxxkmiICG49A0BrQou
VLRWKm1TUGudAYelKKAuZyOL9ECq50nb1WIT+UlpYamNTd+80TR/DouCoyfuuXTwEwvAKT4sFP64
XjOHDtOX8oZ6NIrZCZ+2AL0SNSLWk7/ALz79rJBO0sRySBnfTL121xJiCOOoEtb9h/S16yio+KFT
bTaN8YjWmGUjlrLbCgJp9V9JldMcTD8ZmqWXAB4xOcWHNMl1fhFQaGKIrQT+xR0BxkU3rmvyS2WJ
JvR+dCkyWQB9aPrfdX/t9p2VMyiiBwHshfMUZA3dA4WKyQqn/kGKRqRRI/X1kgFN1jotjlJHBHVf
gunybTED7OfaL8uScaQsRnGut3WfV7tYFMmF4sr6Qc5OkxHfGacX0YCrcpj6vanMa83lfO+72RHY
MxjNLBYKl4Ks0h84wEM4UJLgi5PoEDAEF9Hz09gcw7xzCXJ4a1fc6fwzJ8jITGtNY2taquulHv6e
OE/SbQiGjwYGYnervskHNQfgu789iEM/cjM3mT282xYzswRccxblFSM+93srznyNOhzipjkK1Kvn
JniUUJTjWJmzhAhsuLD8awkJ6qt0rbboNvKL1Eov8UpToxxmvMWzBvILgP+mQzdrYsHugQI6oNec
we5qxb2Lhpo4nw7deMj9pbjsMpInqHTz+zlmWe3F7WzQX0iDcHH0hvZwgyPV+UiBzHk9ptekarpJ
+96vT84m4CrQ//tcIDmviV7bpk+B7I3sGiF+5spN/V4RFzdlt2HeWZCsUSFg2JC5xLJekWZFcuQf
yTrlEsBC2CcgpAH1I7OIL0bKcJacpd6pRjF2UyO1a4KN7jENuU9Z7Zh7vLbJk1VBiXCrbpDvQ7Q+
9NMMNKyRDovV3r9WX+tIUMNZPk4UzWqAuXacJN9t/OYqJfH2ot2PhHbA6U8pNX68+2glbvyRBY//
aB5K8EnaA89pc/Xr6LA5BzjIvChk7kbXIIEilP+og7kIA2Ui8ZDMV8bcYC6mKV32Cw2KwOsAS7Bf
TXOBlkQM14bNqDIzesxTXxoKm4FBJTlOFs6FMA3a7mXTTWlEMg6Iw7JNP5vABrqBUSuYQx+IboL8
lXOM0S1Wmpdy+Cmwc5wN3vRgKMM2t1OHjeiCoFHI9vY1lPJzl1wOXy8S5ydE0Ni82YC9am8NBvVc
zXRNWx6RFQ9o3TuW+/JFJuKR46dvRzM56cSbOcRpo/pHTjLAq33tgnqEOBqhaj6hihqLFysDXuYi
0FvZQigrj5Riuqs2kPO5Pg6Egx0rURFL94swkXQDlBIQK9UiIAsm3zihxHmFV7Cl3a4gqd7TWbjT
EaXrUlkKPRUGvEfaC88FUQCwiAmfyTmp/cif0ELlT698W2MFUfGYqFNDHgeXCoU49ngEMu32Bp96
T8xoWbV7/golvOFle9db9umYsrzJfcj2lizVnn3nNF3MqkWxPzgrID6ki53nB0xpZn/sWAJg4tHl
LOaqp0hEBzbB0NIZ6uOCc5qcDaWeOZJhHxKQyesKboVLr9qEXyadfudxQOBPF0vWMkpXDebbWOB+
UBP7HXiJme86p9Y7I5b9QMZxRM746UOYrZoJWR4KfcN5s/HB2NVuLfqU8qZNtjnFm+W6zaLepUO+
wG63RGiPvAUW+qUEVpBJ/r0CUrUR7YAGRhnx6bgGRi+QXtpDKW7smWdCl6ay+oD+XvB0A1f2Y0lX
W9Ekh5h1uWq5CwP+EeRmGW+Y6f6AGwPv/TyK/4Wq59NyVt9juIemlrs3g9NpOiFn06sgncIBDCjh
C0Jiu8OZAg/9geEGz9/Li3ATrAcKaPCcCbDlauRyuQeTpP7LS0KIeNTWf7gggEoMJ+0ef1cEd7S2
TPE99zUMQvvyWUYVHFKI+H8qSC9zh6lW99RrMXEuWVugd90kdEIJG53SLzaOJE/A3Ji4te78hOU0
/JUbR4Un3+8VVwzIOFVVsyVZel27dbF5Kughj1UIzQ87FNZ7/p4BxzfzDYKSjE04YJBcZY67Syye
0cyzYLrfhmdzPsog5ksbbKbIPcKZXYoPAd0U4h+BqSJSquGGTT8TIXoeJo0XyyLbSRqUM5DWT8xH
B3V/1uufIa84N7GOiIBm1gDx9hLZ+UprqQ6xBr8mxopLAgSBNQQSEKdYIexfqCiYyC5pZr5IQNs/
RDqT5YQBpKM4wyGxeysZgI0x2EWsZr81EEPFDPz8qlYJ0rChAg6ZrhhpVkEIJzYjlC38HBhBTYom
GE0c+E71eIN1tJXZJSgrOlxQFdOdv0Se8CIAFjoSNCKLTeXLkfbO5ITgq+xy13GyImLRbAKd0cLn
HQJLeACL9b6tlghzL5GHyg5055p/qU6mG8aBuzm3oapvVGO6wNbd85uymqeNFLbb4UcpmrWCoQIv
2s1QpfFA4ZqJbl+pRc2O2h1wyQBN6Bwg9keq1E0ub2RL7cIQzYvnGNFF8psQE+wiEBiSgAmWo0iQ
yW3FUhHIcGbk40WP11JLlSR9Rpdkwx4hK2sMtEreJXVmnUIPk/0c0aaSGZtCqMSE73m3rrWZW2el
OXGVR/l8lkcmJP5Vu3VD/ffp2zJJX9w+UpMR4ft9ANq6ci1+/8EJ1y+3iztr1WYN4qTs7JQgOsxD
XDMpncDRBrjyHFo2M/0W/qcaBA4JHn/P6sLwyl0IvfqjsDcZ3HQGvuyRZSinghsJ0DaGoBjodxM5
D6L87VAvpqWrVhtGikNkY1h+kpjKiwP+yfP0lemofyeMMhW5qlzX6vDDLtLmhikLYBSyrOTX8QrE
J+tS8yREZu8vMSK5/gAzhsRLDhzoXF5mlHQCmf8afX/nKRaarrydHAzbWmGHl5EVC4qCQa3lc7jG
w/gbSkavpMVnBYlkS06guT3b8ycghhSEQPXjy/+D9L1arCkK+niZ4xP+zlX9nhrSqlaFq9u+O3Td
m57fMK1ve9HogCW/cuIw39T3GkcMHxLojjzLuCUMq1xBafyIVpu69s9TZIlkcUBoZwNl9tWz3BmP
yuUCkq1rBWqrPOBmMvDfCiVRIgXuAcV4xAWTdzlo3V4/isdn1N3JCTrk1lk/rlc+WMKkaTBJWWF4
DP1oTmosp2g1sYGEjPCWAZh0+n05vvtka6TWgJhl7sg/98c5hF4uwtz2beFpKiu3T+biaU4COtjJ
n4mA/GPKkUq8Ya45Txx+ldfYyJ8m/NrT+hxmvTnom8tDT7vyraIKTtPiMS+HOoqFfy8fuGP9K1Gh
qij4wu22ML5ZIPM2HRHpbHbiGy+mgGVlIDEvyziaqYp4HBEM2S9Voz3yNrh0HU3fri30ZSItJfxK
EqH9xXwNTNC+EFWVu6zXCdcIl2UXVfaBlF9jEPWHdrBdV7GtpS70w4huAzeycMlCebNzn7GoVUqE
oVxBDQyEJmpYxxdYYCkP66uelK3jwCRUxAwN4YW97S4LcKlYeJvQajDrZxpSES1SbgvRt4IlmQpY
zt0OqY8HkOC+Qke2vOvbksaTu6xriI9pbb8eRUzBcyhp3RM6OlLp5G6UIBsLO1XUJteKjsavpdXA
51wAYvUrFcTtgc1p0kT5KLArtjqaU5VpViqQ4IwDwUTneUTTS34gdqXKBqNBvCMg8J2UHGDH7qIf
46MQh3DB2r3cjtAK7N+BaZbG+6XspqohRhBjWJxMGUllV5v7XXzTnck34x794jijV9hnwiwO2JWt
vu3VfzccR86BG/1OV/PX3UdyRdugr63Ir9pmJOIz9F2Chry2QgIHO2xSd1434judUQ16KCZAVFRk
papVL2zpTrMd2OcYww7wcBfycZo5kvK8PR7Ny3cAS7OUnrxQaeFkiE5SOaVRJPAFKp1TN/yQt5UQ
UIIl2pr8ffyccfF6qBwO/EX7AalLV5ScU4aoPzIq+ndNqfH9mO6nlMbZInaFg+F1IGE/yamk+U8s
znDc5h3kpI2433wqV5EFASbSe/zsbs+g7GtQr49C7Y79FbA+dXT2lA4Wsp4wmTspg2uqvpcyjtRQ
TtF3k5yqv/9iqitw3pqqWdfGI576UskkuYk5GEpogYfCh9zvblvyy5lkx5WWwCzs2XLMjm8jpfT5
O0HO9mLQmPxNmfKG0uKrkrCMA6Ad6T7ytYU8B40n/ns+iD6fKfKOGHs1STfkMRkVk9uYpoYYqrns
J4CFMNSGvtVj9T7+dj9eM7QPSPcMDR2F0dsQC+Pj2nY0lMtZ0xf2X8Y8trFXg+ApbuAHKe5yO8kQ
JFv7SqCe79qkWbbuTwXrpuengkem9ruMzG7J3SkTMWAMuZYol1hRAUKqdKMNXRAwz8L4jhpPvaUz
ymhvyBq4cQPXI/2602BSjgKu4odDLFF+T4fqzPI5qjQcAkJk+NZb95X6Tm2muNO1rrxdnkSsSI51
6XKyIwRStZUX9EkBUO++msmi6YNUBihUYxjKBE1uyU+ObCqkE6U6sTGJaP2cfxqPM9KN+lAF4TH3
haSMvILGF3SiEheGlAuCKNDSlg8JUnii7P3GK5Ol/MFeFmotJ0jLlUzUYK5KgWe0MjRjVG0Ejvbl
3Bg0jziadTyTGNemi4BhaHiWirnl27At5Y9jrYlY5rKWAcVW4tCBFR5U2G+a9WFoGNECaohPMPfA
6a2ebxbuVpzYrZpD64VJIT07oKwfyw4RcjvATO2seggSHpniWzXyaEq/ITW3+Q3fhgkr03+QGqAA
S6J+4k/LU205DW4gLhCM9SBNfgUIOsUeISgoWFzywgOJ/Y+ado4CbNsJYw8T4VXDOU3vl9GTPFVe
D8MkFf8ThL1OmG0ggdWcC5e6cHl5cq9Lt5a9kgh8g6DTX/5tt8KvQYA/CJL2qMw0eUgYWvA7hB5B
5RKW8Dat8sgVbG6HdchEH5LIguGpX4pjv01eiWgJC80DGxtZ4P7jMZQfuz11YD25EbJkjNjjCy9k
C4JKxG1nd6n1rWc5LJ2w4oDb/xB4sd4Wi/zOhpXNHWVYhqjlBn+913E2J7GTXHO8lpOKEQlL7xGO
DwC1dFgtgx35y0wtQAvWM8qUGgoGU7FlB6RLMc6B/jk9NeWw56FUxEcxHm23e0z1vJvlLzbHJBCG
kVtBkJQoVurjj0Vb4q7TDofOL7R+hTVw5IKAE8OJgOa+hDTlpVFpJxTw9AwBID4chzf7LMdbFoF4
PtWkfMQrNyX94RQM6/JHxIrmNdKhcS2cQOdkFOEtdCZnLGJFHlUG4iW3WxCSmQYW2FZr3Lda3r0W
m7EI8IwxxLGEJRHDc+DD1WbRcIH3EpGl+lg5Omp0Evr0pAMne/bnxB6lW2yqSJjyRLq5injPR3Nn
gyCPfKSN7nFtFWJNnArFPBic0CUyQxIOZ6AbuCXAAjrhgI/POuIy2WVI6lzVdwXt6h+UDQV1Y9zO
j7J7h1ofdeiSf4v3yz8pAbEURE/hs+V4UPhhjFB3uSAja6EHKAD1WCW7eTChHm7W+QVK7NpiUYZb
yGtJQGeOPnumGaDzx4LeochXIbckujcThPyZzJwb2cfKD0gIvxbmGc3aVZ0+ryWlbGc0O/whQyUK
rYjZRl5nK9dXfCWNLYomtCrkKewODNFpcIYV8seKy6ZjQ6PeddIIlL7wHdLjBcUXUtQxSTDKaxb/
F6wA9L6yCESkgs8W44M7Rv/VBsuMaWoFO5AlXv989Z4JhXPZr1RFQMGEgD8oGk64qMijf5OWObSw
x5rbYf8s3Z0m7Bm/wTWsrbx1O/5ZFoKDrJ1f6HJLs1gaOG7jbsI8U6pEcaC7NEjwky4ubsfERvR0
MU1NeAHT5wosYUPj8WXRcDgUjebvUtw+nr+Gn+6GPX3b+VnTmlSQIPssGKkgxX8q1/oH3NJRkZto
vKEapQdYDKYb/Bpo57HHZpLb2MHCyOFeHexNj+ht38VWG4YLrI5J0rfeWcZlu+VC4hHMNa4psNQs
OHi4NupTYiufC5PU78Jkhkoo+q72h5MkT57D6gJWSvPidXQxCq24ZQ60CPMbJK5474LwlbfY/YGy
MjO27DTyKDkmsGbkz3FSYBfsvXxpS8DSg2kzej2jz96ZVXKfivtzJMj92+JuY2uIAvW2sYe3/E24
cwg1tYcHyai6VN0vC3nyrpEOzMONbyqH/3EsBFmgpF+M7TwZj1SwpRa37mY1Zqpf/0QP2X4svj7o
Jxoa6Y0bdFKPoHtLyo2A7tD9FaqAE3n+916OSvO9KnZH8Vootx12kWaaUEdpffIcFIIdIBXRmtQX
VkxDeeF5ZclJPYojp4WD1M8t6KzRmAniRrtEU98sE6mCPpgwU+dib0Z5W5ivxNSa7W6rRwCsa1T0
pnFpHPIYMQM4btUzg+9tHOBQlRWnm98s+QLqVp8tmdl5eGB/mpt6HsOMDuARJfxEhDdIlZlHa3Rn
VoK0IG6C2Tw+JyT28BGi57d/bsSzcpAR1IbO76fcCGF6l2FhL7n59GSmetE6eQgilRroD9Oh0mhl
HI6TWQF/yoyB5krx3wAfspL3+QdlysQNIyjJokbEk4+He8Oc1Df+Spsr1p2plsW5y6Vo5m9T4n56
choliHDVrONrdSB6OPFCXawNtGtdIThjKXPCR9HdqXmzIjuEcQYg3f5A8VNwC4aERM4SNXAJggxK
KkKMBIPDWJsLP/WJ2fed1BDGTfasV5G4kKw9vLoO5HEp6WQheDUtuudfZSUlYiaFlY2eMDZL49K1
s6Oz1OuKR4zdCbXjvg1K/KjBiM3a9E13wXnOkJO6csjhxq/mkafHEQF0uqf7r68y+i8SjKLS1WFn
UgYsjFly9TZWi6dyWURX+5j+dVc7oWtyQLo0DntUJ/7P/jMrOKESAh89wxECurrY6twXn/RWt9ZB
7sDiCyL1b84ovdbgabdSnGjsmzRIFM00eLphmu9ITrO6G5PENNup/TqB3+xvqT0R8SRyrwwOADWF
uVqHxBrhP0VFuxAFTIxmq2+yNpQIkWjzazD9cEwA1EL96MQSM4laozzTP8Ha5jcwb2kpBtvNGU10
5cJaSFM+lkDBso2R1/NB0pXViMGhojNME9sBZI2/RosTmmqSTuCd6W5pQbAb6Td7+oBLnurNVIlw
t2TUakP0qfc18KZXMcAPvvsXe1QDDGmOSBjT+4s2Q99o48QtBAmN0J/rZGrR1ctlLKymZ1qbXdeJ
EZIYOp5/1FNQNLBetG/VLiK1bYknrmTS7j21faoMUQ4e2bajCtDUzYsw8YDq5Xtjkx/CY64ZVNE3
Z99hiQhu49UV5yjEi9y3LpNveUn7zWaeoVh/V10WY69dZLhc8iDZP8tJrsmI2ScOr6iax7JsatpI
bzSYv8l+dmxR6wUFx/9rSBHisZhGvHNovJFoPRD4qsC2npKquWvYbp3F8ma7DIBK8ZCsdlF+9zcE
/BjEe8KYRabqcYmr0175UKPgJpJKBg9AohFYUsLKBczyVmZVi/EsynBOr+hVGfpMqAfYEH8aVK4K
YUGIliADIjAPFauEK15lCPGmpAQPk9ORXd5gd+PukwTvBDS/ccR7E2tTDl8SJksTwCSxzhlW4jEt
05XaYg7Mr+vph6fIIo2u6iDkMoyJPhN1Ii95NJEgpix3ofiVGnNhmkKXWlp29uUdKLJ1rZEc7fI4
XfNo8RJ3XcxdmS1iqN55K/se+b036As+YVUiFfrNqwVjTyVryY+p5ln043R7dG/eOgxc6q0hcVnU
Q4oNrvvL5uhZ9Cq63/y0ygJu0MFa+0vLJU+C+g/oaIIeD1XoIDP5Y4JabMRg9ojNOq0BCLfFuD+c
lfBQdPfwxZjm0vuQCs5oS64D6OHmnsDAoCMPZ7tfxwkNhZNvlWSI4rlamxnyCG+UkxcrZO8SRKSA
xAqMihez54tGfOHonlRPMrV+pokuyr5hCyD45/P+MzD9kTBj4coxFK/AEYZbfuAyfuqLRQuCxwOt
qI4tQfyzPQJET10xrL0DjT05N0d51gT6gbl7XaPuLfpuPJRNXKCrfCianpAfuBMyoulk4cSm3rSG
12BO/tBEcmZPTABpPf84Eg1962oiLZAI8+cYESaJP25srGvoGUs2NWhVBUnWUKlUeFtxCUS84GHx
TtYmF7KBL8p1CGNv5TUH8D9PE+NFDLNhijAP6g4l6h08pxsXpKcSBPJ+Rg8R2GgEYzQJFR4TIbHi
KCfJ+jDTjin3gMoOvA3vXzk79FiDCSq3VT5JLQvpLB3avs+MrsLT4Ylbqame+nrLOE/lXYwgv5R3
C2tZtDOOPtPEiUHq0nl++xpJNMZSKWpdLPKwxk7yCeTvlR64z0HhfEzch9lOg3yQTjf7LMu5pygQ
Kh2kyjcTe5dgT55drZtt+1JDqgArqVamNGAzByRcBBkT+SW96k4ERL8gOlI8pvYoE1yriAyKwGFE
ptD7X+vr7RwcjdPnrQxdLOW3UqD7qvOkxxDiZdPGUMdXCcJZc3XDFwwMdg2KOlCBtRzddebvKOU6
0h3YIRvPsm7wsdkfd/U7IeeubYIQSlC51PkJm9kITli3Kt2F2+DLs9deG+Da48Px+NJ5bk78OcE+
/ZF4ROD4FdENszEDvVlD1R6/hT2AkfeuSL4FlFzVZsgwssovqm+cnU2G/Z8Zgs2Ee5iQ4RgKZP0O
V6twzpzzMDwrhjc5+6gnLTwhJ/nN2wn5OnZtg6ROL6jEhJxfbGeS+sJLyyRwryc0QN8UOYJXip11
3iG68KUmFDHDBtwzcUquqBO95udiVzuvkz9/5sRgS/yKXizQ5fqNdloOIY35maPT1rC1O+EhIt2V
pw+oQZs3haxIWFVW2l5LMq5ZlvGZZptpe6tvh3ByW1VG1cC+IBY8FFcOosCNeyI2jXbtucboAAjZ
Wh+/CFgtAJhzJCxVXIiD8rQqXJ656W2sg+kIKHZkFzNeAx289+fSskzcYXiAb5Kbook0DOggzMpI
wJi7rRmTRHx7X+qLRGrSyuiuqydhUgc3iMESk6ngOEUq64i8Z6BOv7wiKFClZu7aePCD0uVWDQYs
oplKMoJ0wOoCZ+tTim1O5toeIOyq2VU5agSpuUk+HUVZRzt+rxCz7mL5KT/GVwt4aN44dnKi8elV
spYpEbxECFsbMeXYviEHK55nkHE552RtCV7/LKWMRJQI/VLuqsUmQoJSgNP1wrqG0cmhACkOthjN
Whb9+w+lZ5ZWCv2Bq2DU9IOihv6mw3kgA78eUo6lU8bXuaCdRzjPqfQ0O7TU2Q4I3Sjb62HVuz4W
KPlSVCpl6dGfRtuI6AnxsDcrU4bwOwsixskCMHcaW+R6v9fHSvucOBvgrRqcatF9tg0lHQ7cbaan
iJKM1e3Wye+HBqFVQoLSHyH98+cR4ewgRxSbBUKImEzqKHG8T05Rntpy4cQ/kh7ylS6bfWOSj92f
khDvIt26vwFXyuBn12EVgx8LwHKx+FpJKQVGhaCbvdwq3wseD8638NOUzozYuw8b+UmHYDq3JR5z
dDgHC6x2D+im6xyLab6MbuR6kpZRpzW07RDcTG4yO9czLjRckNpzQK9YglHUpiJl4hBJtn8y+fEB
Ahtt3UvRIw/dgmyxnJHqzwXwphEGYkO7VA9pVhtBqVS6PqDZElQ5p089waad24IhTFnGkyOCK3DI
v7IE8GYWmtWBLQcTtw+pQ6jjkjhbcX7+gYvVlCfV1OH+4OGXMakdG+kDDONPk2azosDw3ECPjRwS
Cz20a9IziKvVTA9XuN84CKSCXiLe44tkC37hlbw8mZ6zNdwif/HuyzuOggHxoYigdnkndx9Qq4L4
qLTpBX465MGkwFvsirCoX3QGqeN3ZA9LQEBC3W5eqAK+NL8aASy8CRdOuyw8FP6tkqCQtQu42fdD
bUTVVzMvcz5kh5buM0nDa/jx1yGVmLWAZIAXx6aQiOTfXpGNAqLKVssuhzsxm6focPiueE/jiF+8
Bb9ZpirGs5qukWpq6lL74z9ccjskR19v9kFXyXjE9AEYhon6lkpZ2vyzW6RKsFW1Jl09QE9qaWIo
hDFRqT+0ArQwMlcP1TJY5IJSNOBJCDMG/mPWFVSVQ1V7B4CHZzWQuBUisZbiblnCUL84qsdVZqDt
Q7VijvA6upDGTgmfR7ZuiE4s8TKs19W48YZpwxX81cVN0GnXH28WXwz8JzK+l+d9SIOXVsCSx+hK
9sEowBdMG8y3U25Tfks05u7y3NTey/RN0QPI9OUFUeoBYLSHOBixx4ZyuYlHfxZ7Wtm1lH5RXuDB
3/eNW687OHArDM67Ujn+tU8xqCOtkThp9UiJZkd2WYyF4fo2S0SLkxNPENHZtbQg1BRo3lIXpbQf
fEvOaqOeWlePSDQJmHOwIy3qCjgraDTPXUR5hWwEg9xMSMu0TH+evvltHzrfat6j6wU0wQoomK5f
XY2xIpXvJKXc4PnUxRSfLkJ+3qmKu7OppVvPngalm1Am+ivBy8huEi+vesot+d+pZOHBF5wDgfvx
lcmoCe8oKnyHZf2U3vRKjYFTqSiRQRtC/+F1/W67zdvcr5qfZpOQlUtOIIOf+9tplHMRveUXzcfA
rtnE1ZYN9fpBKAgRUOsRvpStVhRlBLP/KdBD06YbL3NTsszLJFzqBoH+h0yY5lPhuzu9e8REqZlZ
ywrb5MA83uWXPd3UF2TX65pHRL98kdttRb4Q6O2vfuC/mEj9O+qcD3RZaZWyNaU1NmupoPa3M1Lr
PI1lb3qpnLDJeM0tF0ZbCJl2rkk3m0UzG8rb9mq/XWxsNt4HbIMeX97IDE9XzKSS/V2Fr5RfDRoM
gw0ZgE/jWKTz+TA3oYyaEJtPPAAE2pRQGs4o4EJVLrcbkWXLO5rrlFmAEdb8vULIofoW4EiYxRGr
xhsOBbjIO71U6uxGw6U8hgooJzAorvjlxZVXJUkvlIFigvoSODskXI09QQoNqyp6lieJxiCJHAAm
lbRrtG9rnIGhlqQucEykOPyo15uMYR9781NlnQEY4yyF+cFzMnJxbikerI0fs8ErYQ370I6XgSM/
ELOINDgMcRdl26NqMcQDxV6xrSOLgP57rHyL6tOtzLIEVrSTY2BPT3P+SQhms9dSgqm7UExi3dgX
pg9jiyAoWt/Dd/zJQJ+NBYbxRKRg1ZOeypCAkwGV36+Gr3NL+2qgUuzfMDTkFrzI//OBfld+Ljl4
gkggOW6+IlcLBotQ18bSODx7GFyHsVru9wX0rl5HvkekBNTzIokoD6b62qp4LIFbh7RyqBDIW0P+
ZsFnTsnWVkuhwrk+ozyxxVL0UsqUadSPTeS54uPMG3od28JknOtwAhDUhzT3X/Xv1BC9zaiE4GYy
JvEfQpK3Qrx2/MN18pr9iVJqiGqbrR4UOruJzR/PeQeuQhwSX8rCH8d/NHYl5BMgOBeEdkYI35ZF
DDoowBZ5/+8tgv1Q9Sg5G/hPyVQf/TSxG0BYoFI/JFH773QFWyAvk3RkmSozrvVampOFJwSbCkMM
u2Lu5fbvpWaJEjQTuGjrdtfgoHQch4gGEGuI+Dwck73YpGRTIKpgZH5TlY5yIVaeoutjr3cF00pL
ltdPgD1DyEb9TDMQmCXd9NXwcotrTaKApv29SYxK8equyX72YID2rD+H8Z3BDL1nCNlvahppjuPq
rrIZfJyFoiN238camZ39KSV35fMFZruutzhlkHoYb1lx/pMoxMOgWkxefKiSA4Tf/FHkQjPsmiKJ
wcOCF7DDSUFGkrmPJYR9AVDsY6djoe4NakdG5B2Y38B4SiKjF+yZwdPzbwcp2yFdMcQuaiAMJBLT
JGUockM9Rk8bpbYLmu+vvNYnW8KEF5cPkdrD3qbzl7Z0rvC/tQtWOyaa474sgkouwY4RCpsQRb3O
G5cUA75K2xQWg4xugxqUrSmULE205l5EqpIrOTyPspNWCHfvnrP7MlI1BpC95uNwwHlrSnNvgX3e
tgxp2M219bvMuHLjK/Pm5het1JS9y1709PLbDBFXYW+TJQaJvABMcm+L+pWJ7rmVb5wVnt9GAwbV
5mLt02tB9y1p9MJwxDIeMerw10zDGPZe6UBCR8dMsRo/2g8bs76NkPPeNaErbFQio6OqIFmzJODk
QUaLIpmXHNJER+YeM/il4ZAX6xzRktOIe3r43P+JVnAJ0KtQ89ZF+hqDkQFUf+r54fiDzl6vSDvL
8smQ0mG0y2COq46Z/XLHdqTLXyJo1GZ0bdXNT9BOrAy6gRvlu/0jsacB5tCk7QTTHjdh1zKzMyRH
3YWb5Al+Jlx69I9gbAIkoRmLPCONqfQkhnl7aLCo9biRr/U6yGM3XAuA2Yq2MrrLfKAwi+Brr+st
CC0wQzTi5m4XlAEIhhIVbDNLXKNBFm6uecSotcJNwlmdPAftJMHjDXc1/hye8m6SDAAfdy8zyxk7
+Zax8xe4y2W8GIVuy0ItZdzWcelkQQkWTa01nlnBgcGJ6wFyYOdkze+wDaOjnjNRZZfK8ySa1WrK
daLbrSTFfNq+3lq3TJCib9zYOOG2fem4JXHi9AoGbiVLA5pMiOHumsucNkehaazrE96BsmVOQGCV
8dfHdhVm4pDKWfUaH0Ah+jcsVb+y7pWROG2p7KD/biKhNRbk4Cb1bHyEx1rSR6INbK12bJUSkYIY
eJ53cJLeJk/ndaSuqvKmSUbVs9EJacMNKN6FI3BnCUwD1ubgW9U4an2XW7QeJyasrgpStIq7Uoki
Y0/KczH5ccrW0h+ZgodeecPHAykaQP+QlUei+63fEwFQI7n10jWaEW6xcNWtolm5bZpg/NLHAFKu
rA4tix2dL2dOu+axvVFoIWoW55y6XpOlhyyDaeg7/F/fLWDiq85UIJ/dzu0U0G4C/OvmuHTCvER6
BS6SDbdgf+X9+kbnhCtpbQkbd082rKP47u1zCfuHk8HFQzj4lcBIHpcXHJcbO8F8TeHHsfM+oW/w
n7xniPq21yIJEtdtsrY6FdjXtJZNmJSux+0shaDFpncmDPGGih2L2IjOoV1+YV38IRB+uZGYFUmV
Zrds1YPyOmDKtPr4h/b8ReRWTBu7DjB+5J3Sg9aTKXroXKA9b5l1PE8W+MjMhxmGNME2+6G9Nh33
y+08VavfZbI9BE9M+HscmVpjYqNfaQXJMSGSKxtiu3uH7DU1in+lpqAC60OdKxIQyblW6ir2Eh/C
q2+bkCtET0fDlNC7WWOr5L4TmEntqlKiCfatz+4tuSkBn8O/2NDzNNUVL6HMjEQly4wlE4u5ySJi
jiCfxKqLiCyG+ZP1i/V/ZNhDrXhW6yBuaIhf4WJVBzt64xMYO8/YZe71YUEVsEvOlMnhvw3EddJ2
ht4bCsNOG9c9P3YUIY1LokUqgPqjZZMEccAHRMwDuFYKtSHksGV1s5TTSAp1VlZZvoRqzU2lZHtU
BorogU5wkaJH3IR8Dr3PcC++8m8ADu5s1g0jHtOejzWc4oH+lPupF6wC8FPkiecWIcJ7d/nm/ubO
gp7Csr/jIJIXWBJJl31kMNxO5ng3r1OPHOM+He5V35cPDA2HtPJRmc4b4296ZltrbcBEf/Y+Dh8h
K8Q7SxQclQHwY4n/YHYYnrgyJqs7QOk2TZ8VxaSOYx0N/x/8/DqGgEIFUtnK/fnBtsNOVBrEbATQ
psO9Rr7VZcPFx/JTbwkJTBiPXo/Sb3Z0OodNOZNRfXM5NA6eow8xTayHc7WNFsCXmsZaX4A3sJWR
8xf8jRd0Z+umoq8O3KrZfosYYhqeaE5MNmnFPhRhN4tpwAM0X4LExn8EN855M8ijJ0XZCcSc+yIt
1hXo1g3pexKctvt6d+Nuts7U5vx4WFD5io3dySPcuXv9sLFYT7fcLucNMTPSKP/yh+xhiljX9AgG
OvorGo0kZjG92T4FvEKwetkqnUgqztk3ippvODNn7mwq1pH6eWGcWwTW20Hqq/4+YPxTHcds1zxx
hm3IFL3PwqTMdcofgL8QapEb0WEvCWoLc+jny5SY6oOKLEYqRl2xXEfnlLSg2ZbO3Va8Y1AtissB
fY7PKFksqJ5+ywmbHNzfc6BXWRXcLjVk8IBj6u2aag2otTE5IyPJDNFsuMXB5FbqL4cMkwGxbM1h
OLSS1Lm6e3OVzadLYUVs7QYHYSA3jK3J1QQuaVqHMZUHhqj7s0V4LeXcayOKnmvx9JdEo3mLfpaF
FE/GThUSDt4Vc5Uvm3nZNajyxOC7VhpZ6YbZHki9Lknu5DR2T50YSMhUUgYUBAJJZkzKqcE7UHT2
inAXQZ1wwQ/hzWbuxoxv6KhYVv8NxGZ7efc+mNBvSBM7gE5YHG4yT/tWENImJo1MxYWMrlfoENZv
WV5hln/Wkf7+sAuYxW1nFK0NbofqMyNrgQroYDA9GhgV5hua2dpVC4vX11PnwCjsL6nYKdo5gv7X
DLFTEs/Z7a8oF1KNy147SCS1e4OTez4o8re+fRh8I8cqKf6O5icozaEzZfiXbRUb6c1+8b1xn1G7
fDo1ghILbQsIp1TVCEbX2TtGT87vkpgGE4n3yOgfzVQKpSCN4B3kmkpygSe5P++y7afZazAfgCDu
MDcfKihAyG+akjocKwb4haVCWqn2uEp0jzmX+6rvEmebhscRXklj/V7AS8ku/9QGLESFG6poheLs
RSeHTHsAVTHq1HUYB5VZqrQ4iPCezCHW0c5RrChbbHBE4l8B79UDu3J7T2Clqp594dXP/3O2opW0
PKJ+CgmU3Tzw+VQa2HKe/uMPZ+8meYCb7joxgJ4BQFd5P/3AnU3hhwjHTkzpJBC0w8wDG7iqtYh6
KR9CBmSw2vA7SZAA0FQGv/scGbLmIo4rCrx5GWhcuHlP14pYJ/ZdqZAkQpS+OdCpHc8dZVNsiziw
v1SZW8m4T+TMzEPIWFTl4zgnUMAPtg7fSLWFc2mitDw2qvX6xLsTpcAtD15iG6sSExUBfUbuyTRo
IYNy3K5nh955NnoppPJkknIneWVZuVqcunS41VbmmewVJh2xtca34d2TpW8kUjf5N7Zwmg74bAR4
SstBlRDM8dOPd2m6glr7O4lR0q0o5OcXQKtrUUFr9xEOyTA+COGUu6vGo+C6+DYUp22O5SV38mfZ
Blclg/Z1wfPKNn20GuOTyTH7wfk8lGt0JEUjPswDbMDgAg2ST8/8eCeodPGkGUws3yo6fdxuwg5i
YvRNtdsUkYRgxdFX4/JrzYXWYg432XR9q7tN5CfgLL9AZJ1gwvSPRl5TiCH4Fax1lzDO8jjL3HuX
sV+nv2I4kqy5P5LFAYAOho5E2h/7K5NqykZdZhqKBK9E6QJ0MojsOTro/DU8uaEGviRtn8HKuD7m
MTVTt9/AMjubVjwSssrWUTM6qQvm4aZSvwoiQpPk0nQU43vMe9M4wsWxPbbEHUFMXQcp0wpxFuoR
kkdbMvN4wz0zbuHetlqsN4+nVgroU/qLLQBh094m5Modog+gMrj/uLuqoXp3Obt9wYrqc55hztL1
rOarq9tsUVJG7dhxOryCC02dyMWKGmdJEMlVmLMbeakqnWAiq2yrfv/u29iiBsmAOYHnaOQ23YFc
W+RC40rUc7084Fi5Y6GJzz2aKVDQ9KBzti7V/rf9w4CnCTi1k9XLwrcyojXhiePKhTBA+7xfou6p
x5+NLjyFtkzXDd7INTu4UnkeQp4gD9kpOKJ8LhhPeB/fUkfeOY5duKv8Rw9lY4mrJsBVBs2++8/+
khcVDSA5dZSj0uhepHlTTd/YuQjOvQ10pOynEqJC/RK6P4YzEai7xDafTEacBtXUIPYzt4iZIjnj
GGy27Xgke5zP3iyfSX3wkpo6yZTpPEhaelRNMNfXzFkAiKJiFXROGnid3kjrrLV5eoZUyJPW5/B1
UdnK0Bsh0xDF5GYNBV9IPtaO8oNEWNlXCmBQs8unH4gu8MftANfYr6afbmwvxFF4N827fpiX6BUl
kKV4y8Y1ZZmqtAqn99ccBhwR8dHl3zrJxu/56lOMSKpypQqDVLjCq2xfwlWRuFKb8j/HZGfQM40b
idOJoNmYoYuUC32L82EyVN9NSyD1pQNORVII2A20u7MzOFPWNn1QtsnGLOwRfObQsCmyOdxovxA+
hO5DgGJ4jIfMg9JTpVZIWVUFPZEP4ScR3J2ko4MvVHXhcPpGQW6ExhiA/K/f4lV9+26xNrctT0WE
kC30yTuIlHVI359YMdIv5M3zjuQIQYGaUqfvwsWrbRn2ZbrwjJWU3NsVRfSh6RsQgheVPOjbMNCD
gH33yAOe1YLqw4wNxClSlP3hJzE5rwSTL6lAPq89hVgzoE9ToDC2H1lC1Wdz3+buIaipZnWuVuvp
NOO71hHRYLY7ENQJQtazQ37634XC7HF1vriLw+RebJ+rrDlxvvoDfYWpMQlsJAJSI1YPfmAYdRZn
bqFSp+/GZMRyw9c+sDxvWBcff5i1frLkKoEWzFjEQuHSra69VY5pTxbL+V0ZzYlEgqJ0wIYZ83Ra
sPTS23uN4ywT5YLJHOqHcCstCRuofZZ5R+jY6fF2/YpzIfJFB+yaR/sUKrlrZheCTYCBtczzbLNa
zWJlak7YhVbHvGylXllWN8sB1MKYjmPeAxgyML8Qou0vyMciSQbrU8BP6VR1ZjAYx77W2xGFW1gM
4pNeAtiS6lQ7aiDgfnelV1q81WI2Xe6qwhAMezKlctJVPkitDAhCoiTaesREW1czO5YfsZg+OQ9O
fd9r9leIL1Q8TUIusQ1fsxyTtPaMgpuiJs0wC+mQpy4oYpCESvknZOXqgoLGPHc/T8AK6ECc5sUa
9Pzl4V3OPheKCb6SljLvrF4KIDhTvLfQrI0fSR7H/jdNvztTuGLPLQHvXYHd2ZPIPAhvTyxMHM6j
jfKVJYVccCO7c7NaqnKjHTpZBv+UnIjeJktdeeJQTRaWFKVeSB5aKIRJnhtanXwtcFgF7FHY0avL
TNO9Lar4NxFcEjGnNdxZHZW+r9kSO31X+27CUJLoL8hgejNoPZlxWnALirb2DjVNE9jawz7DliIf
37eU1BjDolgAGSdcZzC0UZJIYQojLc3zT2SrxF2aEULk6XQxvEzS3Cp3mA1qLiEXO87JdKb0chol
qFgSRnmfWv381yd+Ji9l5w6+We7YTXYTPhE16IhcDWRIgNrnCyIyPfoRgWAPgBkRDbasn+NADxlB
iO9DCDfwHfWbwm2TLf0OmXhWLWNnKphVGqni9+EVor7GidfYLokRVcmImV+Cv+bRIBBe/+GoDEYP
AhPkc9aP296QXuthDg6bXGCFP0ldAGLbMckPjMICJJtxr5n/DgG8zZnC8qgBGVNU08k4WZ8HR5/2
L+LcZUyxNBrGw3k9ANp3r4anNvIZxZn0pRAHzpXp+87XKn9gI8EXtfHfobMLmuauk/tECdrDFIez
C68ltGR4SYLV5gbXggrU08KH4m8o9YX3eN+nRahsrJX4xr+KW648yBoK8ucifO4Q1h+qq6VVU48a
cQDaYg7HFwYTav2sNrSFW/HhXiI6OEO/gIW9qZUzJmgKjXkIzz38cH2wLPsxkNV/eCGw2xP7mLKJ
XgjGbnLaawhDVDAblJccml9mCtzhF2UBF5GNV2OOEcf/bAvUH8SlimWZquKH4S2xmPAiHUXfj4cs
fRcN+f7pNrvNDCPfpNYU03/cDOxcaeNHukd96A7rw9Q/F9c8PfWl56llrhVCATTqqKQ2eO3hfUK2
5KWzpTxmk+mkigrglzluUw4uqL0SDN40Fkx6Z7hVgtXLCObRjtahosAQpzQ+4h9fPX4x9L8ndeea
tZyHycmek8GC1qWsSiTFSuy9C1SydEUSXVUtolh4su3P8q7/NNXQRGhlBooKjDDfsMSWyJbHjRrO
pGEd2JqetJW3/aTNykRQsbjLkieTvVPcFae/uXs07/IPDx72d1OK+X6m1imhQR8w/QhxDc7/XAPA
Kvz3tyDVDi4fNbBHRUmG9s8KQgiCpiKetI5EoUxCA02xedzvOyMft3LEjASFjCjl8x9AEFZ9p3CA
0IITIxOVdRGryOz1CgUb9HV0krKNDG29YmNA5DWL/SAH00XfSSvywn+Gj5zLTTC34QHT1Md8md4u
zKjKKimdpj1UXH9CvRNrRPTUhWxiBX5P0nfMnrOg6qU/XdzAFeccsxrJVRP57sJ9LtiTwxPDMzdu
7yIeO5gmdn0qwp0cQY2UGL8a/fl7n4iMM1qhw+Y9f4Gba9icrZLgk63VPIZm46jlKdAFDnTHbx4h
UC+lmad0RcsohffR/ihlUlYgXoDkXK4/YXyLMRLBgJFM5DIYa/81CjGezjfdA6dJvL+VJ6EmdYr+
JOnbJ77WKbEXGD+NGI0UbT7vQNvswwo2W1VBGNUYG2gH/A54ziic67WQa4DSTPwkTy9kLznRH0JX
91075JuEhCGsGZXROE5c2hkBYCSfqzdj/nzT81GYxq2XXZ3/WdeIZJ7XWvACGB/T145U67MHCjXG
PaBhl55gD2IyYfuQWGYwb9AE03mEVBH3jtDe49vc3uY1WAZv6rjpi7h0tFVTGZcbHXAil0Nj5y9+
pTKbqOkc0Er9HWGjfmXTgKNjLTVXi9Nu1hD96x4JKv7VrSku+nlXZH8DXl9A9p5YKg/dAqHTMzHj
gm1cjckJasgLSIclekwhs0vp9L82+ZXQtaa29cf1TFCnAM49u303w69oCDXWmmH4u1TGN5FenKyN
5iB0OZ2qQsmwL+J9V3u0il3Vskquw+dGl/J1WNXFS1eeepMXOB559/EQ5r5KoHiJNZwgF3wuptdw
y5eTmgaGwKhfXjhtcbz4k4Sg0X0I4p7atLl3y9XVwAKcwXrkkuUim/mth932Us2tscdxqS5DV5/G
kBeo7up9K4FUH3XGvkxcFviZGxUeV7D5/cbTezDeQCVnaKBKJBiKJJU6oDInQ8lut+XehAvdYpBn
sDI556EPmy438ZrqjCsbJfNswjfRlhH3/TbVda4BnGLnMj2zrcA4ZXMq+ZQ3RLSiT8Yj3eznesOd
Eij6HhD2f5Jz0QHK12bKrVqwZKYj8MDkHjPxvodLB6F90davCrXh5fQUmIRYUu8CZPVt3imsQxw1
M609FVPoRRFmgIoG5cG56c+rUOgy4DntzOex9gyJRHpc7jLP0/g7PG9SJKfMWXxxsRousiDAw474
Pxhp3+C/qn0oY6DkABDYcjTNBL4aL2Yvag5/q2SGYnUj0oVageeUjZjX62F7CxdsEWiEC5y13W7d
7nBqkZgNBxzt41uRKdVy3wyr7hErivDknzvA7Su3F7WmhDxr792mB3KUzu2XrA62O0OOW2vhcESz
rKy/lntpgWrcAoE7Xw9KaxaglOf3osS2IYIfHSv1DohmoqSxNxPFqYqjiuTcKDohxosLgpKKlS6A
oXw/E7DwD9R1pojszZkrMNblz0SiX1BQa1lyv+Xc4PQ5epgIcW7eIxFb673hwC7Vx0wouzfaFMlR
lNuU+ziW4Bh4CXEk8ZZsSOMok6XpiERfqYfkUuwfjxG39RrsRenu7ZOZygBI0Cr/adxM153rzqps
CeEJ3ON6UgFu4QIDkynSYhtsEkuLtyJ2sLJh6oZdHXhSAuKMe1R8XF3iN7jy4wzLxORRd5glDbgh
VYzAg/ELCpAOAIEuXpS7AxGZY5B3mLJsexNNyj2DTDnPbfJWsCyZZRgXmuYL2jwsoqFqEGO76mrv
ESleblHKDYDy5rGlP0qioq0CPkDQkHzsMiXIHH5/CVy+dfiDg8fWd8MnR0UBJdrkyks/7cC4VEpn
wg1TPUed1KbXtV8pH7bWqTMnQ2LnTC4Q1Ky98YKBpdvRcroG8d2L5Tw7N4RVAqiHvpxsn/874ZAJ
1/Xl96BjadBCrG9PNFT3J6U4rbVqyU+PYMpRjrzUJI2+OrH+5xChaU/34dO7mcgZpE8AtaWkRCJF
nT5uTS4HfYxlFwUtSFno5W05M+CKV8a3Rs7cv63RPQOrMjFsiJZjQHFdfJAZK+a5NtD7IuSUWxf2
oJW/7gRolaQLSDj5I7JG3fjkKHx/J/3GuUYbHRfAXg37mkRkuZMmKkd7JULVBxqDZAXcPZW4Zywx
8mnP1v9bCaHDuyPEzrmhPOJ4Zc/gh+NSN6uDQaiUu87z8S9cfR7smNQhSH9Czyz5KMmJ6/ihA3sJ
eoEe6PVBuYUbdxdjURTIZwW7l8jJOqZfAzJxdUseK1LASzTZiIiG9NeoeIGM4BcoWRDzVo5z03+T
sMPx9tSWvcpdoxomzyWtJo9ZJO8phmxYRUOjHJpno+tf88/5DRHu8CCBtPO0bu9Mc4YXeFVDzTwZ
rIUxirOKCbD9bHANgX7GV/09jyVeUgJWIiEZ1N/GkcU/BLhTRQ+dQf6XYP4IvOIdEpLNlvmBIKgo
uOVNfaLV60ciXatU4OCD4y8lNByAFYM+2QretoCs7tZK84+g+0XYqtCzDnBKvvRwJSbPku60ynqq
/MmJHZcy+tynDrb5+0ZwznEWIbNM8E7F240oqmXPcF3tELTU3TMxKo1oc3JEJKklo2c6TEIfJqmx
8pR49AGqF5WjaJYEIUQQr2CJV1IRmIuGflZuae2C2gF9TKQ6EX0+/bVYuXdyUZhc7eX0B/xLZ5EZ
X1OY5IxpIe5T0gMFp0ugrwbIJTQSDhT5j7ax4iMcBg2ClAMSaww09PHdZfn8mXHphdnqaZQZiiml
JZD8pV/D4NCvp025On/lAsSFzveYL6hHbeLC4HmAQjUb33D4WkwqQTwzriR7fr+xqLCgURdDKpmO
NKKeTv1Qn1mnqCRsh+i0J+FwKIOqLI3IlMcZjG4SKv+kZ/mWTA3srbmQNrLky6fk51wyb2KooMa9
r7c7e2daoLu21tIK6Z66oWgmvtQjkIm4m4PXbfrlbs3LMdXXbjxZjMfa+cGkQVCdIndtzZx+l0mf
bHhudcyMo3xnJIRr3Ux8QafDvP5Mhd/0Ul5GoMXG6e5rirCfutOZsY6HyZ+19uck4QDGOqn2Qe/Y
XIiHLAXTRvGyFtDj1TVZISBejOpCMBp641L15Ne6I4UbR0lYGkwG/RQOGUO9KZjvmHhBooqg1IB2
Q1BaET1GrtHjHhriFZ4vWnLSB9NUO6S5rGksxgiTn/q3FG6xUNaFEtnbOAIh89MeaUjzRLwIbLTE
8dYLaS36Xsc7rDmFZIhhfs5XZlMyYMq6jn96iAf2AMzFFjOsqaI7SSfvIFLaY0Gwatk2ToiaUUYw
lgSyRw1de1AEmiKCTj15oikF0MwJpUW8oRZ0JgUxlJI2eh2qUvtFJUJ5QvqK+xwc4lmTJpjwByF7
dVhjFeITV27m2rDjvKjD+zPT4s0uO5XI/Cptz3P9Yd9Ab1KFnbxIwm7okmXRMont1LsqgEC9zp5O
2f6QZatHJbvlkDPpPU96jeY23CLM0QfvR5nsvQ6KF1uxKJypDqpNcU/QhgGzcLkY2gMY6InKbQ0k
IZCAAu2blY5Tp+7zQvkIiuaYY/Xp7Qtk/RuUo5+uEzVmbj6BMwyXzG7ILwSklyqciNMK4i7fhsf3
G6kfZKWEZflaKf1JuQIaTSzZXUBulfhrW4w9MCKFPfDUwFexSznk4ypiFJIuwrYQaSzYGAgzAv2p
++YCIeUYhznnf5gBoJsawBDTbDehpgCIG3kzLudlnpAfhAGlBnMPC09TPLSv24/1NWyGOvVcqk9D
wSn1nZ34siw7jVqxJWlyoY/23Dx494q5YviKBX9/r3hASjZxZNAyr8yfCoDyumPAq/TeJsRTErjT
fCXfR9IjCLyDSqbCekTtGaXcPwZUlK21BqTO+/4Ssn6uuQGomsReGDhE/LLDR4N+AkgM7DUrwLIG
CAqmsL5m9E+woMvG8rzE8ZMRT+YnUL5zauQcwDQI6uXHU+6dqJ3YEtbRK3k6O65ZKsdSk0WeQBxs
aKWO12flu5d14/i7qSZATA6yRt0COf6bhlKvwbMPJLMoiyVYxRDlHzQkDOTAkATaRGtNYEBHfgbb
NPsy8JUUjwv5zSK6Ab7ogplw439bKlJdmjVFxDRQoTwfhxWgJyDWmJ1ycITXubHY21AziSM8PbRy
z4beU+rDtPxW8tO6jCt0nvBQlUC/rA4Qoy3/3Rn4Hf+wJ+Ir+JGwMhWK4w8PfZyCds6GE6Wh9Sm+
8pmf1lEjOFS8XeX01ofcX5BDHqey6y+ovdAhU6QzgT6DLTc8KfitKHN6EbABWxG9RqSYrBnDJjSI
AZrdvCmOb8uxKangYGqbzcFHzSmt3wKYclt8WNMvT1AQextY0C/Xj3yBWqm7LqGNKPsIW3nw0LFY
zRmOBLWKgs4RB+jj96vOg9PEeJbtHlLjUOZMLqaTcIc92tie4UV9qnum0s95640GFNMltnE4JgIk
rxayotzjE3oDANCx3PWh0o88XOa+6VH0RBTD4lmii/4qSDNJtb9sf8WtztkkuWk5Bq/oOOIRuZSn
u41LBS/Rzye7ZT55qseCzVPigUEMXgEUHzU6KkPR9JDycT/zBVEdy+v6l6bnLNeYdBandSNlXzuv
kAfa7SHh1FIi1VuDDAIjvDrtz2zVx2G9lvPfCFA35DZe5BbKz0YzTa7ncAL7wl4dtR4oCvy2BfqQ
ZY6r/CpsPoCYjr6vmUDz3hdOboBt0mmWlzL8Mj+qBQhKKrxQrUZSB63iUPoNDAHi3+fis5kYlV08
OM755FSgMF1+sE1+E67guK849JDCpnBVlxbgsHHLOC/erfGfhdgeNHAq7cfFcit4ctjYnnJqSDPZ
tKQpjbj5t7SIMWI30bKPzcXzhi+Wkk5gtN6yz6ucR6Dg6lPhRtuMEA0kdN5SQ3hzCifbEriHpmrF
++j0gjZwdvhaZNHThfUwyyBcJTsnO7EBnXPg0TIFLt+gsoyMSwUeUl/G+QsOZH/fJZF2cM8QneYM
CzdnI7dhdmd0al3R8S0mEFlE4QGmeN1X1RH7jlInfZUsEDKqCf20j0MiTGyfwSzKue5z6SIVkxjg
fh4eSyr99uy4yVf5d38lfhVolB/7tnPp53DmxCkTqX/rG0v8VzIDBOkgVNztRSUCD/MzEI/aXEAD
luVE3UhpIU23hpXQv9ZBcbfZdSoqlK7xf8NN5fE8pCPBMa4tQf4WtsOAE5kfmcXpHof1020rr5sB
KPXXbMhgCU/uuTFxNnT7o3mI0OttNAjcDW625q9nFnqyNdoy1dlAeOnVwmgQKKQcdzvTdpphR8Ig
gPzIjvEv4FhH9YpUY+0VrE7P7vAS4Na7mSL63qqz4saiv4f61/4iwl+zYJQl/AlzoEoig/0m3o4b
sObeX416yKY1MkzWVv57IFTzvlnKh/SYDuC5SZBGL02SGzP7f5OF8SWRcb93xFOyaGgKGFzSKHxd
9uAqEzIEh6mCrFngSXfX5YYp90ozr+jUfLJbqgUh8Kn93pLMc+xl4D4d3y26thbbzfJS72+5aPgS
E/pf/vHpRL5KhXhyvgK2Gv8ChKZ9ZCOsJb8Oxq4CrD4+iGwyR//EN28korYkDmfKUciPJoWQXLnn
Z6QBcUUcsOcHtNgJSXXWJp+dx4U8dH1UEJE5fyqYwlgfA+KYMftu8Cx9qKj8S5WhmmlRRkrExS4/
MJSZzFMEXITd2/vmxrMBc21/FM+GFxZ8mIccxcGichjP4eMwBUdL0PPWjaCCcrdtOWw9ipTRfHSr
6ykPR8n23jtB817o12vtg7YMZJVDmP7zVJqXSaCzqiXcidTpyA1VtfM3Ap/h87E3x7DuQaZwGloG
5yIfZUKyqBJOI8nOJGsaR7gYbDfWllktZwpbkiBB84VDPFlf/R/1Z2WLz9by8+NeQnQgGrD8M5Dm
yw9V8SK6cYoCBLGRNUEvHIBTkWhlj4S2Y96gEaFmsl+YatQMQ+Yjteg0w1LKpK8e2AMann6LRbTb
A7e+2ZaM9drct5GFLIqz8sO9+zyz8QWIQiBB4xyq5LvMSd3beN3UP7jRDgCg040iCkb8lkTBmZHn
5cxcTvZwVRGDSedhnJHtiLxUt/P1fvIrjOKJ6Vx/ghJaj1qBSnNmK0frUt4EHm5cm9WdrKWL/xKO
eTSnTIq9XF3bVgheNytroRtr00JFPWC2EGEjqOzMqR9XE7RYn+JBUcppd5YgvxL6B/CVvXu4Dx+z
oyVcpnXgCiygQIXR69gDRwqtDcYU/+AWFXAMkbnIuGOJ+wZG3mAmQLp3smV4j7iNJrOOa3r4UOHB
wLeb+LejQFWCkdf/Y+IZpP4IWpCk3ClbVIzEYM4rcnr4n6e9K/HiQpry+WyfziJ4KpEam67jNVvf
I0DpY+idRFg9e7N96Wpj7qRZxXLJYfT1GNELwpLHVPeDHpRhPEnG1v/9V25PfVIGDYF/v6sQglGT
EY9uc0SI9sImSe33Yq5lx2DQ9LmfbsPC398Mtfv7YVXbXp/hyc0QQkdPrP389pORvVRIczDUzx+5
rXnatpF59Q/8DeUn1N78GEwPVhIZ4Me7BTBpjBv5yddeNO+wILawZyPpJXaka42Ij/iHTfauMwvR
zRHdMJExtonNKdQGCp2uHYqtxQ4u+AecZziQMlNnZN8x6VEAZpbWn2F1mimpQtBAlbT+RPTkYikn
5GXRrOe2+lZ5IqZ/xcFTLCNZjt7QPm0oZzDm4bYw1ZfrleMgVv7vSb94bc5cqvp46uJZy+9PNjDB
acGx69QTvg/KkrslpvhQfpaycI8Tgnn/UdsY+Fz04aY8I2sfdsGXAmClIQjIxN8pns+AgViMd+lJ
71GsLeZMMhf+knVaCnOR792K+9vpGW4M1H7ok1zBT9AlmyI3k0q4Z4i5FM6ol4SCPLG8Zg4OeJI7
ZAeJr8gArGHe6WGaNs4bgcljYaSsswqJZqWm2maMgdMoghelApXrUfwtHWBUi4+QJIuZjO0d63Lu
A06mBWnhgTKaWUOWE/H613fGCkeAnvBcdioubCLdTS+rhIFZc60vpumBtnDqAM20HtnedhjRZSX0
hICZz2R+u+0YD+qAL0HjbbmaGWD2Rka6rWMkgKpXojjp1VkvXsUW9+FPhsOCnrWxh72FiRWIA4YJ
I+LTqZaa52EQH7MMkED5Oszkmh5Abr6uCCDkxo6e3MYOC8I1bsuXWsCIR1AGUAFoqzOYA2PYqJSn
b5JCQLLOp/d3xG1ucr8Ouyh6rNfVjows3/nI6Snv4oOhfl1b8UZFKdxiKoe27Pptq8ownj9WNnSt
7iTaqWp8AfKUIadYxTBkD6B1t1I7W236Z8lm+FNrLWfj3zlymCH/lBPs3U53L/VpxrB72sm3sklx
5YqH2sM1KD397HYRg2AgQejD/tbnYcztaNKrh6mcrVxNdiLoWOfTUp8OcRilK0dbu3V59bRG8kiH
s2Sxv2g3Nx2Ej6MOP6wwtIDME1dhp09J0Ms7TcnkgqOnh5yYI0MlmWI4psaz9Miex+WvsATuJsNO
/Z04LYyYrKVTtmoQsdNyT0qOn0b6c2GvG54L9ZqYKkAt3y19PnRTnAvVujsLtmLOBl+mHetQTQqG
Owdo3w+3wox9VW2QA4w8LBX9XdFvRheyPmE40O7F2u9QPqfW1WOA7di8EqMLgZfQR+B9Y9ukKBUk
6N3SKcwUsCLLa61hbwfYBv0c1R+atT4o2h/lyKuXfZHW7nY8r8DguUHBftCedaWIqpWyoH1yvUBY
VDu6cwag+Hwt6OGlxFkczwWo0accZR5kSAwKZcLhNFKflqndxMW/gLou6ZQzrEFqAzb5IDoy0TR5
/nNPrlNNNdNlLIWAMR/Mv14usoqIV48m97HdVaT7qDxHBMjINphF1pjgh6+ZSuF84bOlMILWHU/r
7h0ygHUKyivckkydtNjM5+WILCx6pkB6e7gSQoqQW/L9eOEQpCo9fw4ExlvWHKPCUzflEvLn+m29
fU6hyUqqmumhWpZNrw8j7JnIIGEzDx7b3zgpaWESMimlZbKQt3ird+ZCWZ88GgIjMTZBcdRhxIeI
SHGMIe1Nkp4AhfQf87Rv0RzA0WK8qTRhfS/hx4rqSZOiJUKyJAAf/dB31ZvVFeZn/hMMkn2OUMlS
qvr2vcSnE/VWOTNc+XJpriVJk+mcS2v51Xvz+FLCauYTuNvfxbvnBJYVJq91zTigBUARx0FUYnPB
DAY1eaUnOcGakX4QKcQ1Ob6JfzqnqPgYXaGNvhVEMmUCEHzI/4DHgFE2GmiTWLl/qlBV9gfnJspm
PiFcwF6rYA10OBf4e0pFy6lM1wrZaPNM8FqKS97OU5tCVQ5BN6QCal0RC+uTc9HijGk7oArZ56M0
LJmSBQvNDu3uF36beTvPOWc4q2hzQnI1dq/JicTb2zKvNMX0rAnEU97v+3NDluNStQi9k+Sf5Hr7
agvRf1MJqZfDsqAYTmprb0Qqqq9tvbiLy6COcvMWHuc4pcmV+XSRVoJpB8+tEt7ZEPBGadIMyIai
zLWRys5Q4ZHS+uCXtShGX9PLOD3jYKvFiCAdcBWTuiD0bRfzGikEZntzyZ9pBztf0wtk49e5J0FG
UH4WcjGeN+l9qPANvD6nq1euPDNSyuhfPk6ck0/kq/bZf/ajNusDZT6btGWz5mDY3KSs430ZHh5p
NBWOUdsAHm8/0VGa6isbpRXJa83qo8+4C0Gr1ElQAVaykNRJuEQaU4lW9uVXssl9m/SoIfgq27os
rYTNwU+dOO9xw6befeg7XRiPy4rB1+aj8491vxGFjIJh26fnp4UuptkY0H2e7y2Y6qvgTMNch1JD
7drWY0s8d1zO8dTJn5X/8XPnZGhnCA/c+DdZfM3uj3Cp1VOYAvtNT92bEaY2q4HScQ4nV7XH65w6
vvZ8K8m7iC8Lz290ChsSzYDp/cws6L6otEx/GDLfBL2qozK07Fgjj1SWuZDmQwNqDfd1t+TktmNN
d0OL534CHSKmK5rynRxs9Tj/9CkQzmZQGSq8NkXepzfoutlACKNU+AnBKm6eNTWkObQQobez6QTA
EZuSL5UOZBprJ//PL3y8YwpdDS56mk3Y9jWxchyFS47lm5021M1WPY+8ZxPK5sx04sLPJaAP+MzL
6BRNDMSjkc/1t+BrYSfcITN6UhO2OalmCBKYmDcbFNOkIG15flzukGScJf9ukaWNebmrEo8YfYjg
nCvK27rrKgElkV5pEikZrHwLayEKJvoRHOLP++8mTXCLskShicgLP1S8DPlZyC76mk7pIGBwYd+u
0M2dJzfDHtrGyw598eWVEYwbhwqnoKqRuEMkA9XN/8z7y22bm4dUn7zAzZkBMhwU3sLZTB7KQ1qK
VS4+8Qa6YE25pIod1zVVmlfK8x1D9Lc7r1vuPcvzZHiJ1IslTjDaPuXmtb7W95vWxhKtFuZVAnsd
j+Mr0MaZ76AOMtV5LRWea529fjHWh8QdM+AcuiF+CTe7n/sdoheZoijBM35roPnVpWbkEBrYqlMZ
bqEU0k+qZdmfT4M+Zuy71jA0M7G9hGqsHGXI1/CLrltMs9Ne2sfdGs2/8XK0z4gBN4fJbOPaVIa1
+DilJwRYuHMaAMrMWuTJBaBd1AYBnFYMWiEHjmKtkqrypudce8D6ejYfAGzBbLzKO/Ea5R7pmMcL
ZFYw5Z3p05gv4moVmu/HYev/CFDVdmbceF7z+Uj7vbRUoLb06/lXp3q7FujRH7pVZ1/xkPJekYZn
q/u0CEwwSxDjoeM7aTe79ipXFM1Xt0sHtZXppUaq3uj+b00OaV/pqZZ9IfRLPB2ItWNOCZpj6vHV
M1taROBNTLVTQHXk7GDcSf2LBaiIMBOunYM6OL6L6ziWWl+YEgz3CXTmQfpEUIBbIVFGyOUM9xyX
P5Gl3ulL0FBZSaPDwtu7b54I6CUoEEUcS/paaLrIET6U4eYg8P3435xTyYP5rSrfg8WvdBV6mPEP
l32HN9AEvfZJP0bctvw+tWX3pRh2yONiERPkRGV6BXFWe9atH3v9Ro3F166IDQAcS/8tuvxTD2VN
YRstyh8ZQWdDXS77riW7ifCg3s4c69xpKBmBqH0eQHDq++shlUoGCdr6iogqeXNqY2gRdv1ipMC1
X8mI8QpSrSh0xBXXwjCVv+5qxJIRdIyf5SOZmsT18nBPg35n8GaWIovRb67pyw0xk7cWN40INTAs
Fr3FrhYTz4UPSRKvlrSq2DyE+vxPydRiTilkAqwabh16SBLV1XHTfaBRvxQbwAIHG0mUW+iWwJeO
TYiDPYitjlwltNEyfCS2uFZaf0QdvrQ1zcr0x4RJ8JK98qqc4et4MgKbup7feia9/s1MIf0up2vA
hc+JhkCecSiaBLX1KA6+iQUo+bvsEL6ZHQ6RhSH8adGxEUpPDUtWUWtbFSXJTEZ+sGnpZgRRx4Yq
FTfawl+0pseAeG8ELlcpWeh3roqR4iYDYYLE8HlWK2O4nOYa+tBcJX8szLIuLs0guii2Gg/aZ7XX
nk3KwoOE+/Gu4D4eSezcPlBIRyyxath1RExQzmMxATp+iTRBKERF8H6CM38I55ArgMkMHai/nSQe
YVMM1qJXTly+n7JZYyS8c0wOkSjBWz+V/5KsRIlKVxJIduyj7nPa4OHzVHYuxi2CYNKP2lVlhiCq
cYEplUPrJROazaOcn4UqxtYtFrinqehKfG+V0bNvKHlBFhzSKr+/Eox3/tiTR5cLJrJjUlEV2LkQ
N+NESvlGUAinu7yyYGE+E0ic0DEJRCJadwEDDQYxKNMSM6yTVoFA0LCmf/GFWD4jHcVbRVhd6Ldb
4dCWEvCY95UXoi9hshw1mx08bJAgsTTi0NpXpi+7B1KRwNs/ZriX1kkE15n1z9qkIg4kX/nJpPUi
xNJ1RBPGZqGUeQk+0i7o7rR6Y/iCxTVRTRu/PQw1m+CTwCob0NQvD1RtKkUKumSEtAAZ1nKY6SnC
wHwXJr7I/iWwOjm2LLCoHNVS7EuN7VqY+qdHEGPYEMxlfsnftG7Sj3yneYm3Z3x76ZNT4EZEiD2f
NPsUdLwKv/HPgm4gYeYCbMdUzj+xR+QHF4xVeSPB0ilt9rxq6GyfBdELFMoeP145HJ5zgeJQ6Cck
sTLJ4WaB5QHZZom27U/PcMfEM+u4bbn/CEpsGwtgZP3XNKBLzVxOmsaRR7LqxX247qkmZZXqVR/o
/abCw0YWIJQFGvpJ7N2mWHKWkQIwGTKY5kR5yM87zgVrV6zR8ivRqXQRFXN7mw71Gq1NCe4XHJ2o
LqUQiN9f88WwGh+WrHk5xnS3XE2m65/zIqlo3TOukJDgMKVvu50gkRwWt0tS1oXObV0kZjLHxTfb
MhrtROyIx1CoZTwVULAJLc9XyII21Uyik57zCB7WScxtmua/UwmKr9a8REzn9Q6uWVFRDFJTXF71
XnLusK+N/UAF8noLQgfwvjVn4yuybi4zax/odUAkwr7Vj40DDn37iqGqve+rI8GLsTY2JDKlZgFf
1vSD3bPVSPJFawnKkejaIIxIcgD3TpfrYJ/rv9TATDb9+5oxtd5IuNTH/zdKERMaheuofTGW2Bez
in5Wggw2Qma0ScXMZ8Tv0uDMb0GwlBgii260GgYv4uaJzJUxB2eoTM6TvPGn6FFSkYu4nX61kdWM
W2zd6vqGgO1VokQGGtfFhd4Qxv/HOtHxdE91ZGlmio8A3HZpM9zw8aLoZ7vHNcWp2jHwcjga0/On
SFd42g7UJMIupgkTmGbiXYs7tPM4rGIHdF3rM3TK3Brua1spkSm+tbFWI7QfoSVZqfV2Nknz/nni
fF+M3worHr3K5/24Xy8UeDHtsSvVMu1iD4My0M6M5oeZXHtSfBKkxC24RmFGjs7Wnm9qMB4mHF/X
R6PGXRyzj110Wdx5ktkr0EEFvkafqX10jOR7sT3jAmNiw8SUEQyblfpwSUxwV8PxNJU1suDIZIk5
NAIigIH8o89hT8JB6vPhnb3qJLrNvTGOiTMjT56zWsKumRi/OS6qCfDDdNcX3fWFgEq+0tziVVzl
loX0ehkCwDwUig9oPNllDWGdGqBBmC8KrMb/2neGoN8FthMPth+/4GwqTJ5vvXAr8Mrm/aRJHX0S
G3rRu+k6Jen3VB8oiG4je12CfPBS8auHx2ycmR7ocowna8/NaEKHJ+Nxn2lDTftnnGOdrzE1p/kA
V6GsGjMkKf6fs05cAFbOUoYROSVn3vhP/7TddAI1gmZLl4RQ07yp+na0kcH7sMdB6qow5jha2pUI
e1zHnGjJ+syzOTuH4A78Gs+JvEkjwbxnNcR7D44qTxPdyel/Kr8y1sJXYeAYzWv2Nzd/V01yuSgI
8IWcAaXfjFlhSmuKmvmZdeDXReHKfRAa8uZC1y4KwQn9Mo9lJv1TdvbwzI59pbJiPbxkGWu9qYvZ
FlG/TLcIoFD8/WQy4QHHGpt3Zxd7dSaZnlkbLlBKkbiN21dc0HVmrHIcpgWxVz4jij9f8+ooW0IX
0nbiQrztABWRziG5674cQ8wFb8Zp8LTjfL98PBfZe5FICfiivElzDHLb47ldfKcbhYgCsAbUya9I
h2PiNpZ+l78Pg4iIbRJ8ABQpNPkP0ErjnMxF5svXrMKFVXgJQVPaM3nSdrg2XhYvCjlxE8SbnnY4
Fs5Q0TcEiz0tXaX+mMJNT7vqeRYwgu3rmQA8s45pzMEiq+K+FjkaQLx4x9mjAPsmAK8D5suhkErS
cGPj02+zmg4qnRRiENQl8vcTwQ2e3V9KxZu66TdjNgv/l106THPc980YeoG0nK6v8ielYz4Zc20F
0dKXffwb5XSx/7kzSsWf/JXHf8EnahCUAC5k5nFrRgbLYSRUFjlcb4uZ8OOBoR2586FaxbjK3IBL
AdNZ56oZu3+1ywxLHDH465AwEvEKbxJSRBciuaNu1rQmBqxMp9GiD2d9zocbjr8LQFL02Vj1oZcm
ja2WptRLYgCTp34OhoWks+nEuLqX3CysEDjSm4F4loXx/3pEvsHzhc9tzkWT9ix5IXfVVefTZ+m0
jimMU8N0L9Tk3TXhh5iUrc6mhHVCfFVxGvl2BBsuXICJc47IjRb4YUYhFXwhkKQD1jBXZn6SbrLi
wTddmtg2Fci0z9lx3eeeab1FADq/7FkV3leiVg0xjvGerHRjrD075FjpmZf4YWDFYptzK7Du9C77
kuqoaRzOzTCm6GOqCdtvt/NCtxDe+Meiyt9a09Z4EG+BvgvhNpB3uG7nLYrPLdV71F3IvoRu9hs8
y3dih/VET/dYSQ3sS2M9ztWYd354ifdmvQKZIl7VqvHeKVTS8HtUAl0NYn5nJ9ym6wwfnE7BOekl
j6HYK1iK+uvurqLQ7g296/ojbrlZt/k73eUj0vNvaXxQF1lGHRffB87iVEpEGzp4U4pVv4EBxc6g
etDheRAHy/tauN4nG65qUGzLBYgEMOjP1BLA77obO9/48QiTxoeq4YGgr0Nf3a1VEp9qWuCgQhmM
o+r64Wj3IYeeTH7SxiFkKAsCeZ5/7h39jujKpPHYPuzaG3x7/mpmITr/eAkGDQZXy8rhKG5/08Nw
GSrfNai/8EFqNw9pnPSiufr8sdBwi3sDVWM31WZVf5f+Vr1qeenHyFN31ZoBawRAbPXHx3oYXRqj
C+FC3G1ppGPPcE725bngcNxeceTwFLK2HQbyF7XUqa7NPOQl/iKHo/y8AXmfqYNCVpGZIQ37E3/u
Blig2a/X+vXnP00gASEkXXsseQaDXdBUViu1WF5p0uTVjx3HOsBpiUYJ9i0JTHgDi44wheN5jqon
iIM2J6NXWIoTNMoq13JObsh3G5Khcr+TidK/Dpm8YNNjvOBWb0Q9lazj3YTJ6OMzZb67NcMrJKfR
/C3jLQKB4f6cBhqV/4lm/Ci9BAk4/6k8tBd1C8mjE1Y6xHJ7UE5YO781EZevTO9oHz9lzu9vnTFa
9tc0eI2NtTcKhf95Qw4iV0EOwMgdK+TCAzZe8mKc+e02KTaS36xAL5WO5sZ1Bs/V9hpGZ56/lXCC
ChmjBmMxgWFhA34LoXmlguyfqmwQ7fI9+0DIkC9eK9D3RZTzkAZ1/JUnFS0qIVRUpr4PZSiMQSd/
qGIv7jxnXZEsssyzqwRAvnU8JRkKimJrqgdUWDuhbQaGeAUOkPdLeOWaYKy7nQK6yTl/IOD7y4ik
ISdDEuejEWVxhBRDWhTi4e/Ag4Sw3KwayhpkYNzQGl5rw5LmeEnLfjLqXbYLtyx261hLMmkzhqrR
kyjTS/UF/K4PjRTn7bxYCOnRTBKDpGJFlv3oLPd5UV8427asX4m1UpgVGA3AZFYtDLkX2hoEqf3a
rFFzCBLpIUSmybyy5g3weAON/Id0/V8oMUVqBka0iAWTXgjkFgDJ+TSlG5aY8NLun5Bh4azxeXSA
+O9iynqQd64w96w2czcbocrbUnA9AwH89033D2hvwjgiWzugjFboyqbfu839vP1BHlqclUYrGLOY
efndMePgiQAyZ1zNfnxoZLJM8bjMc9BDJbEJruvTPuJ86zwNvsNCkf2Ft8SWIqr1s6SEcrshzed6
OmHRWlWwkC3WXd/SLbdKE/zd1Wb0YnYpkaF8cV1nbv9g2dKMg/l9mql3MOYJYUeVV1mRXcRuCyfp
7vimGI45FC4On1DmX+oBiawMDXEKZznwMBfTqxeeu9+dJK2VbTYdwYnfKtTMs0CPAmqmgLPBcd+B
czlDyz6SC+xm7AnM5BH4T+NE0Pnv4mnJfCI54N+4pCx70yNxJPIQmffgHf3iIh2r3sJ0Ru1rsd7k
lgHJ2riNoddTnbpQo2sEL0bJNwcMVMSWAzXqZcYQtVFHmHOPl3UmYinOrWOPOG/yk0LxunoOz9BY
z0FwWo+rGMOCPYAEDWbuZH8WSBI8NgyYT7t0gWeqaMEV+muNWHAwcM4nRuK+JLecNGJsZp0a9vd8
0FiLpI+giVXNW2W6kUrSxKj2mBf4rTITZJ/AB94Y6aU7jnJTxdewF3jtSHdVa3kHdU72YvZx2NoN
KxGTRGdMPoBztXO+teNNk3qinWbkm4R1Qk/Z0+mVO8dBE0bB/T0fheI5M2ZuwMsQBstxIcahAWro
9lV0rN7KhfI6aCmoSzeXNWMzQEnBugOMRWpgQ90C4Lux83hVwqFtFNJPr8cK41IjvuUT3FLxguay
2BMdUdVVlaK/6PYoqDdHQkvvaEKqPQU1R6pcz30jLE9MlwkOy8edmrJndlVCDKxkL0TMfK6SnA95
06TxH9ljlM/laHbon959xMV9/VteupKIZdEJynFAweoSHnTC5TpxLdemk7N7TqjdjTY9vx5OBl0p
ZJmGpzTPaQrXobQFUWCGXFR0xjSwnJFRi6/05NZQ3GscpAcPGLcH0fKaeQNyZLTbTWDEygteEX5Z
2zr6w4rfadWF3S3/0uZag5tNsgMLo8fSHEjnDFUH+Po3WVWVXNLtl08qit+ggeqaY2gh9/QPAagt
Qb6skvHgFLv22pm/KaBDHfBaiEwsDfjv7x1RyeY6NTzfj5exL+ZFQ58VY6Aw3Dn/ycUboHFqNQf1
pnu8/Ke9EYNkvJ/ZPWQarFzbBtZMWUIxNF7fGH2hVLBVdCsD1VeCR50U48ubvLWRPr0G1bZ6kKnS
VRdy9tsv+acjlfzvCUP6/kPLsUFut70FSVb2dW3vaf/xmJtMAv2oZuA05Ky8dbejrHHp6H/mIrTp
JB26oVhZx7iDCTMrnk3Q2TrkuPQuR4qrWwUbm0P3MyZiyV3mBalqXqQH8VZAUhdsdnyfBa7d3ftT
1cTMBo4EK6F2apkMC2Z6GZd3VORYnvAu+Q11LEfWDgF9ghPBSO3ht+fS/YydFw0EwvtrwpDamtLd
p9LKu/ifDlrGe+0YbSqInbu2IxlI8Y3FLGybjd2/oIa0u8KnMaaq8ZnHbp61NrDGmI0OXQhLnzU4
H7IpxI84YQzNSisOErutVq+X3LeKyWoDDi4fM8c4hAfLW3vvnBABc/kffgiigSSViT1EdtyNDB1b
2BqO3svKpbA+8oTTn+wdT/YbsYyZUTmZfFNePbxbUIwMMT97E4IL2TjNV4VK9jJcc+ny+lnr1n9Z
NGt9wkEyN82q4rctn+3De3l1z8rHsYOOkw8U0yf5iPLCJEKILH1J3yNDm5JAv9rHnd48YSS/dd7r
8T0sT2OX0becCdSARTOihCldhyUtRFWVpcUl7D4567ZzZhEzVQ2y4GqoryZX9mtzfYSm0ULgoLf3
OSG59xBezsEICUYtFNtpWZIbS7p3bWq108Q2O9DpZRPBs5E6t/sXZzBggK/+O1W2OSS3sRlr/hBR
+S4yJt6gw2IuRY6LeS9niXq66TdqGIehcpAwOXT19ZYO7OtnHYTXCBC2+Rg/uEA1LWpF7ZfvyCdH
YNIx/wpHwvUq4VanJNKOgnIJU6rgvAGAQ3o6/fk7DbdaNFFXJPPmvdZTqkDDqY3fFK0FTg7OtZlu
x3pLJSEBipnLQVCjwTchz1VtFD/W0ugLVd47RQkxJdQsWGNUJEmkuVnA9z5fxuuJpougpFPkCmKt
+tneDcBpqBfPx68UBb+BRfbDljCRESu1BY5WNceQQDUdh27Mzxa4awM8Y3dxXGPzQxaB1fds9Vqn
4c43x22wqUgXUdaECx64zdXNf/R4jsEeNrOB2vtzgPPUBymvUFqAzHH/Vv8KCd8jv1JFmE8SFzQi
31ckzOvaMoFGMh3eBK0sT8uyTEHiXveqv5O35TcpYG404Dlh05okzt6J25LSV2xN7oLdomr2O1wB
ldqV8us2hiZjcaoFlqHPRX9GQjHXCrEOwR/r0liPC7XeI3n8QXU/zpMP7Nu/Ps6YQ2WtRgi4AKBZ
akBpco3VBJQ3xugGdIPMW6B60InJrv+/wxPiCo3mPJxyEwq7mR+8Bh578cwe2ToGYZQrHHfe7454
W8bVdWtSLCrslno2RuqArmjibdvspzvkkVPnAjwD6CAZysVZq4deVNoa+CcTyhODFNad42jVsAq+
v5inI1M2h3mFfsneHsG4WvgnOwhOi5SC3vUvuayOBZmGvGm0PJmuuWySQGCSf1DaopTwQ1L5dEFm
EAZEUEaIi8o7N+121nhdSDLOal9KZKRd0BzEfqvzFqrloMAKWPmn+b5SHFJc7vV3y/SVPGHvJzGA
MSpaMdNpHbZzQCiYjl1mnEw0Vu3ZFX6CAR6HfZWDhpatzG9C8u66KjGTw40rUu/Nu1mx+JOtGYx8
bBc9cbFMWzn25dyPJE2ciZjaBwhw/RxZYuEKkrrT5Z5sHuXG5SVJsf66Xy4QJS8dpcwsV64v+4Yq
2Zm/Z0PWthkIe6hLlMOJErKPCOOJe9rDsiHq6WPw7xcxBG9gE0wbCQx4kkLHheeLYWKKLmOVGCFx
b34VLz5eTUqysmFoF4KKJV2bU0kTGlE4pFEBupJVDO3SZjGMjaM/fWqOqP74n5Cc0puHTnY0NxUm
ybYzGM/TmHq0wDX8QPp11D+jfZfSCKrceX+hP2nJskCK9Q8s0Psk6uuPOx3EV5aYBiD7Se5Q81IR
v31LsJF+OwxjXPoj3QJGLMwiFX/psfOTVwaK9w2nqKlFvQQ2sTg0peT15hIIzY01VSizGI/xJ88e
v4evv3JTJXz9WTMgFe9PxJGPHoXHSZD0S39yz+8UWN9Tgd0FdadB8Y5Xo/4CfnbSzLoZviD4OfhV
6+6B70/xgHyu8NMRX/ZNmcv1NXfrzt4WQG0mzl3A7Q3owNmF1YFz/Eu/0oY6B79AOhsAXW98TUgF
jC/6nC4itvxgV2FfFblWn0+18OGh01VxlV+mZZlzqCsSMZNwBzaoDq7WydD2uR8qFPf8CZGL5v6B
jP0gYIrStrJQ8R2KhVQgvhBGpV2lT0Y6/of+QpKlumGUGBnymgXQIXh9P9NaueN+208bIBQJw2zv
11ORQ5cfIZRkKruVWVYenXECQfPonmwOXXr8/f2lnv/T3pmHcxBicGTmIHcb3ZSY9jAzdGcQuVXz
5rItLswQcSjm4TAfiFqxdOMoDmv3KxdMBQfoJIXwHrGQxUVAkZRU7X1LkaUm7+2Jo+L1hZTgJXO9
ICwNaYmcXvskowG/t7j8Ct41OuYCaqxa3uc/d2vcI4eivovprpf7KnVFOuhvSBolRJwdqOIwCe0H
0EX9Rjd1DlY19UMySjwx1YPIMhE5aGgT60nq+kpKObzFLMgBSQj4AH+UbjejOzGix90VUiEcXgEy
AHz1bpUw8rBvXMLHjAY3b2d6VBr34tbBhmVnbUxlJHeiXpAvad3QgMgh4/a7hoNn7iU7tyrvA87B
RIadm1bwo6a4PsGIx9OwvSkGGX8g5GLajqPICWbJMVyRSrJ2svxQNA3gY9lyfvKG2SOJkafxLygf
7eXutNjd0iQwrOC6koYpSc9V8KfVn9kg4dkd+Sw5qxdeV3eaB3NKwALwXJTkvggdltDmVVWdowqr
JBiubbBSFI7hda5ypq0WuNCssw51slRDEVj909DSNM03FfOgncEZGyYsd12F7INd3pc/6fmMbPIT
O9Lf2u+ZfICY4SPJRui3+Ir5No1VdNdkb/XGLOww2C1KEnufUEIbpEMw/5b8sPFn7GhnZI49NnvR
L4+VzBqj15z4X1R6K+dg1sPZTNtGGSWD1hT+k8Hsqxi2BEzwYqYEEN9tNhY1qbxOiMsSYrB6mgo1
fN2c9VbC/B2QVHxiVB1gwasqtu5FocxuDRaXTPWTurfcB5/uxyY81xTAdUWYUFDgV02RWqLdUqnD
VMhcg0eqGKAbn7u9zjA+2p9nGdfRTSfEFOKlucGer8psGwhIyQ/rQCSSBrn7dD9zOO2G7fZNTIRb
VgNjsfJz3t+R75wVAZpKhoDiYRGqeY21pZtQc2wgvlb1IKv2Ds+YLsaMiIEf22mX1cNwRZ0T2To2
EAtbzaih3Tm+LHjbSNr88p5sOIFih/iGBXMgds3XfVn7PNTE+LRkmzWfX5Vb7m46sP1vRCPB6Th3
6JI5/9QAi+0Ms6vwhcnPKnReJGy7udiorhkXY868tLfkBcCI8DEcW/OuqAKOGxNtZhHogFfr9Otf
q3XAV/w/WiHylvY0ExXpMpMc5YF7Ld4kwRwHHVFDhzS5KPJrgkUmsv/rpTM3pWRDyYYAkS5TJ30T
JJ21EN5nTLa/ZRb/d9XX177Fg73+JM6JEMCdc3R3Go2olRuOZp5tPXLN4w1BtOgE4PIW+0ekzOIt
QONWJE0A2VD6+I2yDPNSM3+tnia5cqjifU5zVClcBpJu3JpigoUpCDXO3U3jZFakEULbwFyG59Dm
VKop3GO9g9U4DdtSJ1bkzcB6h2snqfXISKY3Z7yyLFdikGxC+RgwgVzY5yoQcjAYwYsN3aPepirs
Q8oWWjjZgU6i1v/Kv64ONqo/6zuTBHcp2Z5ebpmZsi3oC9iwgJFNiNV0iVvrdNBVD4HUfPMz8Frn
KmDmoYcCk/yBOZNURpKie3QQCTCor7zrvr2yG2wQ04ldyGd/wBT4qXLVBY/VZfnGwFxaWlpAHRh/
8OHqawBNtmAXmiitdIC9P5pT5E78z70OV2bqvpcbEUt2lkgqKzsDOBHs8kQ+V32ztMf2MsL4qi/F
nEreGx9M2Pay6kVqZQDlUCJMy6wX1f1ONVFXUv03erFmVgmapWmRRLmtXmRlvu/A3H79FrtGnRI7
C76B0KXiOITv0xlciLE9bEsh6zpGk2mvWFx87f3pXJXctBiIogdyir/dTWnMEq1+SOi5ekDFT6jg
oljzaA4sO4fopbqxmnFJTldj346OGPY78zjhu7dgdWX3TGVdQQX8OFEJXsk0au0b3BnYdNggLfgq
e2KYwHcFEgU08uChCv08VwJrO/ZdL7dhmrvbXfWnCIhCrAyJP67oLATHs3bSeCkEi6ys0JHMHYn6
N6QUAYljTTpTsIquJd2XdC+TFPBwo42Rk0kmvghwhCTySkJBAHn0gHF8eJYObg1YqEmvAcbXUPVE
CgnBtwUck1jZKLCzNnuyxtxpNdO5RbvepkvX7t28FO46YA+zya7qmY1k1UyR/y5ePSYMS6+DcQQD
7dIqQipbhJEAcdllE3qiOYktbKQz8DAx2AuhiwW0ep5/AGIR4ozXnHrESOK/UfUP6IcVdousIzoP
Kypscv0kNXkZt8sSu4ybtQOE0fPZRhFDbAx9+7UGz9GMce1N1ya6uBdt/c8W6ChNoPUzRON1OoVR
r+g1UTgP/1J9DzYWwQUOZ/MDR7846H2uyvxrcLOCeZggkjrMWB055Ne0ubGPrtpuZnUEWrxBtghX
qCKm/Q3hHMry4KtjTQXTd580doqlosp+UVGWed08ERtaRwyYxWfiYsFMRg6tcwRKRYhXORydjyx6
dq4OKS0g0I3tYYms11eQO8yHbYvnyGFy1Vn+XO39G8w4axF3MAd8PUb+Bk9K+LIl4P11TaTlZDFa
kgBOssgt/4gaM2JBq04RN4EpPKAXuVcxqLTlSPub+F8BM2haJzxsowmofVZxtT6D0fH1Iss1kFxj
QIXNOmCwuI6NwnE6kCyxzV7FDwyxwc+tWBykSrLL/8aG8Hx+9xykBN2Vov2soc6tJ27Mquv4NA2V
0ywpALcTjDIdwqlPzPEzvUarIbrNMKAS6XxWMJY5Dx8boJrpEp7QolzE10fIZtkOwRyRG6eAnVuB
m61/q9zcgI0bVKxihSUkqvqLs6ZUXTnj01fD2IQ1YoC+sdWIxFx5JFPiwUD/vZafLAIKlTkUjpKd
r4W5ed+ab5ffYvck8yBimXodSZ8iYqlgh2O1KPGq7cSH/MN6SX9pNZOdAB+jyFKnHbChMx4zyczH
o5M5Z5hlW7N4reTzrGkWm98GHlYfaLbic7Pt7oUGKYIQEYAYzF+VTHHwPU7OhLV00Zlq/iuMUXAW
T4SKC9/OUgWkN68HixG8CoklMJPvHmDikLOb+oGbhgjMnUBGVbtVJ0jMDV+De9nlv6zBTY+b+pjn
05Kkl79onu0kjnsvhNVBijLLUB423IydZu2rvR+QDQx6XHwGIV3veIjqTfDUyc1GBrFoU2LJGTZr
sbcA3mNU+XLW06kCW/pbfiDlmvuu6MNrTCrdvMO9pnKV+pX23p3ZwCWW47uxSmGsPhb7gnwwHPrv
/gzB1c0LvMkvVH6CwMGrbKx8k3qAgrZ0udgTVS/KgAISVet3kqFfLWH/L+dt23nyOlyo1rMbvv58
jbFsGRa+88IZ2FUAKdhBw1Jg7vjFCDNV2+GNr2En3T8fSgR4Wmu7wKTqZ3/P4ic4V4pxR6a9Dqa/
yFRXqeXKOKhdUCDzZo1uiitroVY/JwL8ZqgzmIOZ71yvo1g7twVPU1jloqAZpSx1fjXUVoDxNeya
ow+wpXghQQ/V9SGscF2Knfqz39iMPxZhltJr1ciqSNdzeUNs/RopYqowRSoFc+6Jj4NCTTGzKvNV
2VuMzw2/an2GLI6C5zLLGFgvU7WitVnOKL449gIcBiFOZsr2LHZhhTr6zszngKIqyTFnX6Ti/fRD
t4czV3xOJn6KYfa5Bv2er9i/yPh5RgcoB5sPy88eTnP5cYN9XTqXxxShpT/6jSVrMDb+4pmaAH5G
WNm9sXysplqJBQsFsU008UqofPnRRd6BUAS3Xm+RRxrSlYUh1li9HPpavIGL90LUmWutn7nsVaM1
eHAW9KSAGeKwSWmziN2S9fRV5XCFaCSi+uN0BkKV4Rsc5fLgWvuMaXwE2YrxJ/bs31CUK1Wst0EL
3uXwX5BIg0WMrV0gUHjFLllxhz14wiBUkBC/YVF/U//XEUZKJqiQje3XLFPlDfekNjDL6UX1ZQGs
LW3RAql5LH+ObJ9YzjFfDrvyKeUuA11dzyw1o0OvKNm6Mu8ZgMGVAIwazZTY6hW4wHTAFOQQsvAE
ai6i2neBgczY8hZ4qHhvKenkpS830J1JGsdntm5S/JZ1b3CFdSZl1UBPdoAhNx8V/kgWlYegy5Qm
OdBhwLfECPorbW5k/y4FF3orRtAVty9uN0GCkST/AP5AVOWyPKs+NG2hUo3HaebltnujHHPxwLML
kkpNbN0qJxdl9Pc7AUwuZjnaI7taXfgy3dogakSf376+zFJ/CUod+kZashcWbEMZMcbhA7M7EpG5
u20Pdamg1EjKUlF2KJJAwitdHq1YGWFwUFmj2UfnTWpw7UWXFnM2MkH7Lp/DQt8/J0dBiBn7Lhj2
2Lg8WVEAxK70OO4X0VQSHuWDHjsTp0nLTDeQ1t/Y5LLW8fgaLQiIWQn9pxI/K4woRFDiEnU/JNlb
niAcxhuEZikon8lVFCoQpOSmosgiarsqBKNetO8Aqe9X9+YE6DWHC7YVnhGqGXMNow1a91EnSN9R
HqmnWOVgJ2wHyDSRJvdHj3tmNULcpDGmJCMVJa7IrPnY60Kw6ym66qeu7GhZ4zwdt6/jfpPAAOub
jszHSTAOmTYDUSpvUljQMW30qsz4+1MVcQdN8Hyoc8QbveemJT1WbZwDlOJAGKKN0kB8Y75zJO86
eOIr8lLulqH2VuMAcsxNqlgBaT42QasJM4c55e7j9GAUCc0U4dnRU9Fktcen2etfSNYjAcyEtc8u
5C5xF9QpbdT8EwNJQKp5TNRLHHLRb4paMR+LPUsT/wIozuMWmKSUKgeQhsvjLahTuHYoAfmqCxH5
Ak35Chv3kRrK3Z0dTxUjJhs7dgYSkvUhfMPIvJuzBhJv36EVfj2xuaDADge4RYiJcAKtnjfBPbOp
Ym/ve+gucoqCwMMX+0M8csSBkFlEuXRE5h/OBJDRULf9NqY4mG8ssCkIlWMe9tCxoCMFGcZAg8hW
ZZ1eeohPnBVE7LgYBr+jZumaj94rl7qxUsaR0Mj1IL9yItH6bbgkFi0AlX8pM2cD9snAgh46AwB7
4q5FA9WC9kxHSz+5K19/E/RrTQQZ1wuCygdVTq0ammXdNMmebPoX8fzvvVbc9IuM36yvEN+GGGER
kFIcqVRhauS1mKdB3JMYW6TiEhQGuyCSOL2/FN/LHVt+YsMr76pFMXYp/fzV+Ulb5xZ1t++wzEUC
h0gWRbVX1CMBuv3krl0w6FKYJkdpMn0oNXcm/CxdbEOGWYPiT72ZGMLLo/znLZFu5qSyxS2P6WUn
dCAbZ86Igy5FEsPlyt3i1pTrWZX0+lGsHZoeqFsQmlh9Fs22lbpRCeon/iHslS4JVRA2ra5JA/Kr
9qgeGhD65ETc3z0r4DL8xzniNcMwff8JEtRxGNiE7jzwAiFlXDILrDMFpB11XpI/CbVxVg1lu6bl
D0VawZJZI/HGG47NhfPMJ/cT4z0lfFqebVkjKIJ/fcojzkws3fTNv6X0i1RHFwphL9iqO5KGj7g6
hlpkl09n7kTsC6EoT1GFRey+9GfSLfqg0jbtilaiIgeJVLGQX9Ugt9Tqlw35mkZaYWGyGWmP/rCD
vujFD8pEFfe2DIXYGltBMVuv8NLFlDsQXUjRut2tvgUfMecn3MPl3kW74EC6nZ7wYkC97Us6TkjO
QkndKdFzcMdFjVHs8Buj2TAQCEo5uYTXbdnRPcR+YAQTksXV3A+XQ5uc0Yvj0yzqOsut1cEkPNbs
mHqT22H0NP46V5BbLEBedwk9Xf1ETbXK7XrVYKngjkLzb0YgHdZ7NtxVAz1s0n12tG3i5gaQuWeW
xYmAbPrE8T8TLt2OadXfxw8Gh5kMD+tk86HzMKp0F90q1ykb+yMZxtgTbNiP0lglIOzD/w2WCAOP
6GAYsGFB79uKJ7hvb3XwnS4FKTHrfyITLGNN7K9uvSPh87OZWoS1TI0RuAMWO2cIvs9kVSUzO0FC
r1WT/JDhmhpfM9XGzWrHYtPlo+LS2L9u+HH5Sz/fWM8aWiWNPOK68E3tc1agSOlyyQvre/WXOspv
oduF45Mq/jo46gnj/ms92ljEWP0nNQDpUgyVngf2BZvKVIOUVf2KEDzzfY0Ajg+QmIrz5dmofUCd
xInw/t1oBoLUOx9DLJtOeQD18gtb7QyY6IeMSMZ1pdeQVZEhqMDkE0X6wit/fZPBJ/8SRiVCTtSg
3Io1JZLfFkF0+t30kCpbDxR+3rE2sH6SSItQlu+6aDevbDV+/CVINkQtm4nHw0WCSTBjwftP0GZD
0dLXslYhnNKVw5O8jwBowAY3S+7LEKzJT57gEXETzPxLdAcv/8REM6S9CTPD8QjtzNboluYuk87P
5IfCXWP8tTf1/bcNP9z+t+F5eQ7k/f04PAm7xsyStPiXxvaWnjCBMFsDfTnQg42raSPSMXQQXRC2
MujLNGd9nrQda8AjkE+R20vAbdAJYBDUFnRuHB9tMZx9oj89i/A7v6Kx4tpBpM5r88r++8pWEW1d
IGfcU8ayOcyOkfpqXCqcbmzFXXrGrHs+d2ushoLEZg8k6BuL7pE3V81EeGAa17vmv8GQ/1t9rsFI
sBD9/zThSfBfo3vC33xcBeXFithaQC/4/y5Jq49sTxSyffRmMJvINK2D24BP5wPJyDKaO78TjbXY
R1mZNOD0E91a7oXCAw0PeYLRgaCXCCwPpBuu8lWn+eYjibZnqEAW//pG3QJoIKQIQILXI56pMjcR
/S2fxLkYoc9L8qLMVWzyIN/nWM19kq03UYD+S5df09Assw0QOxpwFZ+yjSE0PNdroh9lXXwi8n/d
Tz1QojKyoOHrGJkFr8Z814Xtemf1d7+GYIQBkimj7gISGIGbkdUzwVx463tORPcwCCmanpVs5NN7
zab68aof2jxL+hvs1R78Z28WCguRj4nxUELOFr0MUcGltEq06x1RwEifeiWww+vIJ4aL6HVzJwow
EyJ5USSJGzImDJpg5Yh7jGYIiR1phMrA7teJCKvZxg1eiaj3d1UGLwu3Smb14bKj40WPJ0tUoa8b
FQEh86f0yX1Mjlo004jfuiaq/xEfWZ7SaLvNuPEdeIVGvT2iuWdFMUQOXGYqBs+yojXJnZU/42wG
+soGmuC+MH8p5DQWNzBnJ+ZeR0Z695lUGBYOjIIHbeXhKDViboAC+TqUtjnteheuQOQiSUCjCpVz
vzr2q04WBZiChB9eu2Q+pofX9gtdsQVS8BLcd6+9YWCS10gMcuufocULXfShIQOd/KYpngX8pIfN
2QaowGkY154M5RjsUQaexYqdCCMkP0X3Rg1LMLFMJDUDoERML+2BjMoUrhSbq9ZmLkHFD+VctL1E
tIj0jx/sdwuJGLetSjwKXV7qa7CG2nJGEycBQ4tX8+PxEJwTWKgJfoHvQvwWOKDA9dbKJq5LP4Qt
bTHz3a1VYTRxLoBZsrFCL51YIs02malm4KAIs1AYwnv4UYhq14HJBV7gEjzHOCEUeEJohNMTG9S7
z5jfIkyJOAiwHKZ6UlKKN0IBZW4LqVAlkKuWLwrezRfMDQnk8MGK/2BmOKG9LyWmCT2KTWMpaAKH
AU/a0/oRnU34hBNS5zYa9Vjoec1te0b+UQ5bdbVNcGlvN2aGQzj7Uz9FEDlcYriOMIJ6zns9mWET
WlwcTEXJZiRtmum9IE48oH61AGuuChSkTM8dBU42ndfpzN3QDnkq5qdzFNw+Lum9B/ZzRGxVRlww
cNlf9aHk59GyiaSI717hij5Npx5IoAZMrXe+9iAJlMnlTl7UkXG7Gl9e21yjDp+94yRb6CtmZQTU
hxBEVkP0Z/QtMMTN8nfTVQlJgmQrFko/2yH8BxOcuP9YAPXYdLfKe00pXpX++qj8YevAqH91eWSn
7E41mOQDSuNI0nB+wglvFa86ZmdGzQ63uMdUMzEL4dd6QT1sAO5Mu7Tdtb2brRMAXvmdfdHJKaUn
FKV0Ddc7hQzI2xItY9H+9V5CkakYJNe42q2fIwmbl0TICCyX6F4fGoteyYxuXKAJChr4iiCYTvPl
Zly7pFCUPFU8ZgnkqBcDQPVo3oVnxQJa83/g+tzzJ43LvF5bXgxH1DJ8InbBwDoGD8w9PQqu4bO5
wXMtaeT7j5XJqk0QeuuUKOwXrDHC5ZVayH+1edGaYBTosVMUVgA6Da6Ch/ms9YQqwIk0Yj1dVHdC
cKHsE1VgJr+q+7si/KsoLlazMPGb6YZTTv2FOXqLizha7Iz2PRTRCk6+AqKZX7oaoW8Hq3B13Pa9
yVrWNwmaBTknXLJ9pcB+HA5lC0QzktteRPx2OfA3QHZ63QPY3z5jQXdsjQHZwYzINJeFkWnqCCvf
GUhHTJD3COMV6Og2zQTEtKY1M8SmNSsfkR2vJ+ko0j+DcTqexCI3Pc5biRwRcqwHLnT/fJx1UjXE
NR/vePwTg3anzVzZi3QxSGR9OAKTggkQ9lF8Bln9o0ipmx+/Et+FVTkDOQ2PWmXHYtWnfdkNtp37
T7L0HS6NUGWMTHmmfl/aEPOrrUcemj4CC4HyrTS/8RGo2NRNGLuJ/cwi9bZ9PSK3Oppq5zca/8r3
jhdLmJfKw0vE3/VKOxCFpmOq9HzMXlr0z1BjE2XFzta39mdQtwwxpH76LIGVFthTjQmEUp4Zi+Hs
oG6B8Lj/tMPxjoXjU3NWjZEXdJamgugnkQcjZxY/t8SqbgFomxKxKZ3HFJawBGWC1dZAm9hhbuBJ
Zw4OBPZpyXth0Qz70Ju8DX9F3A3o9yjoA1cYvYgNJkgJiz8QELGZv+PGTauwuCg96cUE9MpL4He2
zX6WILXfdTYOiLSUA43RVmCr++c0NrtB/9Ebfvbk81zUMviC2qd3i4F2Js5M7Ae+P64VdYIzzq5N
M6jKfHsutrr3PMLMH0+VKL+75PRJAbm/ZzXodWN/o85FMFGdPagC9rPfuBIP0VVASjxUN0IxJe9L
pH3DuchAPIDGEYvOosK9SD8Ewyyb64+Kj7ksvIA8AkH3Oi8KqWr7R45NMu0oabxL9HezAUJVNrjn
BGWCmEZ7OhJd4aMHuLPDCZft0JRSot5cOJFda7tEBQRC3/SvQJ0E3RFk5NEnSr0wfmC8V0rt40Um
AfNdXkxmchgN/3u1y9EobKWI5u9FzswcoHRB2ZtKlX/1FLwIKbDiLj2rXOs/qdJK6xCpOaIVtn18
v1LCcAGEtM9gpdV+2QhIvLl7/s+UY/vetrx3EVOlEAbjJppIxYghYZa/R4oW5+V8krAIvhcM7WLP
Gk48XSGcYC0iAK+sZL0R1KdT1ZtwZ4wfrCYYjWH93n+CRTNVHUpvole1Qmm6bJ8o+i+Da0YEc/4j
Rl1lpADLoS4xZLg/BJ4fzNavE2GtQsRePeFOWUTvjSP0gM+ebFteRHaZQWZQQnIni7FPrSMmDLqt
G9iOEJVaBpE4HkoDmCODQsYVvYamkUa88OQStSvmL6d+A6zeQIQYlRM/492EE2WUZwVbuwTL2xka
0qbyEiFRsLRTaAdiJPBtRJ6JRz/KIQfm801wUwbA5l8b6EoH2LaP++exWlrCG0WAzwxWD2uc6HgH
4nPrHKzJo0ViLvwkelH2MmkVJ9DJ2PX4YWBxP6pT9tQ/6zCoECDadrA/vXG0E0e4AQC+GKXeeLAo
NJ2HnOhCXjc/Pk7Q81OEJ/Y0NQX47+WDs+qg9ZAAXzRn8qahh3/u0dPdHZ1eFj7M7vlynI6uDz7C
5QrDBAc4yZVIeC032s9v/nQBAxoCEEd17ip9oTm9DFLenOaIW4rZdu8NWFJtfyPEeEpWaD8itHcs
P1orHTiAnGDHFglwF+zkzI8eaZiHPnEP00dYQNejMWXZLbI3Pu/BEHUIqNX0MDUNXuZfE8IQE85w
ELJQRY4cckmBAOe4zITQUjz7Zm9YYAeEPJYG9BhOAReWvPrGbx5p/IKWzCtclLTskuPVubAt1Z/t
wcyGEDc0oEdxn4fp8mGNfL5GDRupJzEMnzo3yZU8BiotX7NhoI26rNr63cWnfR4PbhoyrZI/3HQb
444H19LVqr6J5CgOfnqgIyXKe+FM70ZM2sjOz9G051Wngqd/rZlBOlHhGRn1Shj/VV3Gt9iyQwm1
+r9cLo58tm4xIvixgneX8FkBABoYtJ1TZbydtu6ERRiG8/kvQ/U1u8WqMOyk4EH/jRA6W+fn6BFa
vcWfc+U1DmDW7bQjzXd0EFN3jpC5QEJJTmcEhAenRTK1G6k8fOsNFuJqL2st7uc4lW5Sw/VndKGN
x3KaA4sqsOdPDzvzEY1IuootbSa4Hx5RWWkorfov3XoEdKnw1q0erj6QEezIUkvW5lsCO8wIyKbx
UABll9gd0C1VW/ME8u4L7pNpsEy4E0MoC//8sC0jtLfEs8psODOYZFWYlhBCYgPrKEiVTM3h1L5G
776dQUSaL9wVdtSJA6Xj3z0f893zfu78NK7XwgKIJErXwYZ585Nnunjwk07Y1KU5fUxBOCgzr0tP
i/RWjwQ2EKnmM85oz33WFADFWJE7ER/h+xO85b36sqJlxTjPFRdvv7qHWiy7lwLzl/kPjx9hTzpt
EPBHo+tcgG3YQc5Z/RB97Su0h8PrcDsbQCVLZZB075f5cHHVmR7ohJB/iupIn7hQKA0Sk0JF29qG
nIDDj3XVcgmYzOUNimq89y2vP+62ZG/I5EKa0sXeUkAK+JMgPq8MF+Tly12s9InBYu+ZJk2+4XvY
YHKtn8jKwZvJeElVHiqAlaeoPhPno9ZUv8MQEOgV4F7jzsflnz4MZ5h8YgucjKH4/3qic5m8mdV9
t/pT8aYPQQFwWn1tPVRR/GTws9NPlFgDAiUpOpPnsaIzQXd7Y6gfsKUa8eLUxoUfGk8vV3+ypiDN
huBBtKn1MOmZkEyjDca0BXQS68jksyAID7gzDi7QQ6TM5OzLcKj1uz8Qa1AK1rG78JMnga9Q1Jys
rZPR5+V9y64rT98M7MFKJi+ACyGgFUTEsmEL+DVBMi4kl+p5DIrO6yx2qCiupfxxNtPmPh/JUnd4
9gIA/9TcFVbSEieWtBiyGffva17aD2lgs4OqGxlQsNmhyR79tIQIHKuVkgCH2+pHBDDs22lcyEU3
yRHswcQdOPTLrBQRFcNu1zRivnCDNrhtbznB03M4cPNEUTb0PjVCQH87Di+d+zkRkTnuODxrwjr/
kjerqb7RKfgwybu8iavm/0rAjqrma0hgErRQ2kLE7oTybWX6WBuAXBSjySZ7wm5cR0i6UTa4tB54
6/2vffzFGdff0iM2BRbCRSuB2ViDks3l0LEUVcAQNst0MDSsqRFnuWPh1Ug1wwIf2moQJtPbU7Hm
R04sI+/eSSBP6RKROPGMNUnX2c7tYvR0oUytXbMhLVUsdpHqppP5rUhkM2hPy5DQdVBybsk761dc
jS83QvQCQMbLFYSF4hDEMy3G2x9pAxSf6G+/ucZ4T67tZmbSPJ6jYqM4RRmxil2DleI3Fjl0y0Mb
wt3VnZ80xEUnkdjtavPqd9nmueT9r8Jtfr61JoUmnIbTMdyEdTIUBlpMNODaWP31W4JKlLLkScs8
+TtKTRVUeutNjrUQ8r9kJVjeAweljh0YX6caSup3+D/pt9DK6/bQ9LfIvDyEhYHEgSewdtNipVNq
pMPAkrOEsplrEgEV+YgtVmXghGhPh2joBo6VlQ/aHRMTka8dORc7RrmmQEqp6OQ4q76Y7HGvpMFb
LWwz59cjag3URdS8Gm9rPYVypj4ZgvnB674t+EIKU/ixgwVaaOuPsdi3P+/2tsqlmhvTG1WdoV9N
pe6dhcuO4lXMoNwCRx9PCm86mjFOc/q1VqVEVrDCWBJV5Gu831rMYf1bhLhl7Ecam6chCYzScEQj
lwxBMtAZleZRIRTDJ1Owf3YXWYFB7AyYEvCJ1OYTVoXr2iyXykJa84YCF4yUkYZwL4UtYBDh0Gn/
ZHOX0UMHzQiCa2fw1Hf/TjnxINgaXpBLRLb9KFWlVp7zaMt10/zLRDTqzqLKDR+lAmYOhThRzZQi
ntEaWbXNLpyB2I0evULvaV7f4KIQ0hN6rY6OtDDSbf8Y0OvZ2Ytt3KLmqICeN//0HsEzTjtmcAC4
P39bNnKV0ludFb08wW9teWdCAkcLc19ueX0EIMYmz/uXvqQoqYixeij81pQEFPPyn3CuGpDnzgAp
kJx2dqWvodCGjOarSIs5lDmk3N0eP8lBq2s+TJoxTloFt33/Ejcfz20XQJ7C5lDM9/vnpvhACkkr
bOjXmWylfTD14XBCYRaCvnqXGnxUbhYtfPH5B2E1rUrJSqs943eRUUb9yk8DXd97DTfS1AAC7uMy
DMqVY2ZK/XLx23yHo4/+A9TFG4kYm7XJOmGp8Xd+yRF6Gg5+iTX+e7A4flYOrK7BZlWV064iMRsu
K5l1UeARAFPdSutk+czyizbGN6lFWXrVRYXYccKC879gR9/OBN7iafDSeTeNZy1W6IkyQpKGaEaE
lvEWkAMO9r2pj7mbbxUuzCPWw+hKWEXC/IrWu18xjsYJdF6Wy8afKXm+l9B6ae9XJZLoEPux3f1P
H2R32ZUlTHkNnQDTGMYb43GTH+s1FokKyPCoNBOPIpgDqrEAi2wC2YFsZBh6yXTfwbv0tuVyjWn/
dp0Tsd+iBeClONA7qgO5iFu79dl1NwVQXTgCphOLY7RekQP1zJixhJxG7RH+Sn6LCNE2+co5HUeg
XBx5rtb1vHlCUHT+lhZlBZM/HSFa0WMn9KAlOAbeSuy0S3K+6SqO+5dg1MyO1TAS84QcPiYV82LK
IaBFUzJtFQOwgjHrz4gTF0C+XTKwY8s4j6osg1d9WBdDCbmlkXtmMdqGdmUwL2YlZWsqEmb9kiT6
ax9dgxZunIWQ33N+OLlQTArQEHOZhRd6GoVQU0/fmSed78LzOsOTgjTV7Mg5dgHDiyP/o6dvo2pf
n0vQbW2DmtQ9ZazGV2HV3b5EqIoLar7bg0I+4hISBJu4EaQ0vK9ttlpdwhNvYxV4fm8d0ZiTKSFq
WeYLz/ENuTULS5oPcBWd+O4O0+Aif3Xj1DZWbRQ1j4pMNtswt/jUYLUB9PAvjxr3KwsQJViFEemp
ZFrUDSInAi7SehxdyimEA0RKHtEAgxsIEbBZJlROyNYi3Xbp/8mIM4KyQ1uXhCH1a4kzt4X+XAkx
cZazVBtSGhbm/9mBIqw+Xw72B5Qnbnb13EzCCUmwLDHCRtUL2442WI6jjkyA1fupGh4iwlaoBovX
2SBPMy8K1t92VbLOYgex+PSMs+dD8tUbL/zig4umEcFUDzKE9rMzxCG+QMiojPe1yMQfL564Gjad
8lHvr3UJWJJTiUjdnn9/W6AY2Xdkke8EUF/TqZHHz3atk06hzPd4BlAsJe2WfuTocHqFIfxSiZu8
HZ5seqn7OgtdjrGxay6sLzKVNvJS1dAeM8R5FcQNEmxhqrcsKOFxniTtkxe82Z8fQRvn9mVHAqeL
ZBtVa+diwCDQzWpn0UqYTc+mu+6o4/WCtiNxRdcPZaFBgqK+D9bdB4OCBBfx2+hrExSYQnA9hZ20
cI8PUOKtIrLL1SCuFzu1LDejifTSGkXUjcf43IsUDBejNbWnlT5Vu7Qp9fbw9UI+6DCSZsR2qzWC
qhT/0LeQe2sKPFKs/LwN1++ZOVjE5B+4MqloHsxGJ1d12AujgdEyaIHZid57PKhaw1lxxUuliLRT
C1jrpqLHqZZpk8X5QSWPUyiemi55KvjZtX/doX37U4yatv8chPPieRkggCpjX30BCDQALOxlcTvN
0pPyWIM+KIqk6GUZvfLGxkLxFM7rQf4Vu9lGBCWTXHiUyEdsGA3dfIaLcFPLyVNqkr1mf4HCWDlZ
xjnIgFPXvAJOP5KUBtau4pttdDY2WGwFXWsFOM3G3XLmY5qg1QpNah31ekeRsbyOTohD/qcvnxQE
WV4L2LqhTPgm3hrogRgZ4NYDG4n6vnb8WaNj3RMTpLW0bdkCNmiGaFp1iF9MTB8JsTHo44s0fwfK
IDZKT4h5WYDQTHnVrVd/jiRc26jJHhLMcVD2sCAFeSX2iN2D9duzEA3feEtRxQqEMx5WTKPL4yog
LIYvsfuuWrT4rL3INDNTwTtzF8OU4o4eZfpDt94mn7g+t06DnQaVltKBoOzTXwD0hpuTIYrFYk77
FDX8pmwBUdI3/uOlwvgnpm39lRRRTs+hxY5M5Cs7yD4Z0wBxUiDZB897qZTKcqcEeXpbwCipCznT
ACdhG07ZXUGgicq2MT5cwNvGw9mmardHSat60oQrVcRZ2NcjhX17vGZB6DhnAExVm/fklzamWQoN
wCSAWBFkRrRS12PS506ey99eAWd+4eR4BiIzJzNJDyupdmGXaZjdi8dFJvRHkfzwCoEd8Itu5l6D
vSOtya7qtlB/D1QDbHgRerYRUf5644xKOR4eaAZ3WQOPFUkM+HuYZK36Q4GdsRmAdw2we7Xnszso
7fO3OeMZefKmCZlpbK/Tp5wINhtaToqsVjlj3ygoVxIT7ARZjr/OjsMNs4fyq3tTGib1XXgjvc3t
9XdF/gQJdYYjEJhaVJm7MHqFiSH5IGEymx6FEjF6dntd9SPrdP0fiolccSJql8UgQfIDTLHaUrul
a67WUd6LIi+rNLk6vGuNoEOSG1kt80PRx7M1TQl8V6gMNkeKRss2NPgn6bVRE2/EKoMT4mGD9+ES
DaBPP7DH5ZLuW82ewF+A59PX33fkA34lKkBxnVHh/2v3H/y891iDx2dSrAbdQKFc1xd6yW8M3Ni1
lTPQMZEIKXxOoR7x/5ARJubcftuukD97KA1uGkH/CSWlFxPZ4zEnRl5pkSLkLGfLlHOiAqLgWB1V
dNkJ66b8t73z/azJZ5a09K/VxUsNnNjMq7alYk4FlkfSWWX87QhtpfaPF7GgqU5kiCYkW+BpIBsD
WxQE/BDTRQSe67amoQ4abvOAb8b39sjltDZgukS6ejgQFlM/uPkpDD5QzYL9gcFb5BodtDESNz2o
t1wWmZY9Ovd/p4xMCWIx6GqCjoslo6VHBaQFHe30kBTwQDInHfStdNgKm8PhOO8RHsNJCUUO9FuZ
xqsGFxyyKDsEh3pMKN2qFFIS1Op6qB+u9PQdmsg8ShGEKEIaDVB0/qWTiXlfayKBAndpirz2yuOD
VswgdLhUFgL/seY0srAyuytYJ+TxQ1N0dVKOFfACP2ol0QJ2Gd4CLICWfaN16eO5n9a7rGb5guBh
8Ic1UvyguhP+OKAW8QDHrecSsj/ROhB9VqLdow4kSP4V8UhBegjRBV/TwItKaCnzeygTgDipN85L
am0xW1yBfYg8pepqpWZqFX5FeYLZFhhDXG17KKsJeO7hR9HAWGMBMB9VfreGVVzYuylpNvjPkXg4
Kzu51/W/uQnHCFxzT1xtfGzwOcs/+ZhFCyIlvXromM7TTwLFgyCaO3lzOLmGIWzduovJqnGY32yN
au1gQRIrVkxupCqRGCNSo8Pne2NrTbqwA6M6diiF8D7YIAeCwJhzZi5tzaT3mqTq72i0cDFnrv1X
9FqmcjFcCLpoQSX6/mI7CdYOJnxRgYE8N1IiebRmqTY0Ip5Cd5HOVJMggiMnwsCsIcyV1Bwhyz3v
aHSb0gnMDHTpRjPLInOgpMRFN0rer6SfcF/NtejPTJt7BCwEfpMzz83FizEkpeE3+T8bS5ijSyCr
u9V/ChvQLgqIA23BKf88Fu9mELL907GhH5X8RGvWtCt3EjQxbZWyqlFqBhqmJSf5ldauhoxKXHYN
kgv7o4lcH7N2ZY33ct0N+H76zMUWjNPPYojT7bsqZRP2wBC0b9F/R8a4XvizqSj5yRRbIVKcDp4c
3fQmpldMuOSbpQPUDjf0qY3Vklm2nUBA16rUcg03TUCM10Xciorq3uGVCYfPT+zeB2DipDMdjeni
wnOtwafH+5YQjNT1yDhT7QiM8TYC1Nyrx47MZvEO4XvfxFavtyh4XK276DxhBrd5bdydHkVT2qTF
V+U7Kbf4x0/aAEr3jN6qZ5HKrOoicrNCP1WyUM3poKEGpRE5+X25mdKM7E5FNld301VZH6WW4Vl2
eGTQsrYSGxRQ0h/2629sXomaofFsNaA91BaE4B+vAtyNAp6D/Qt2aWAD3khiz2NL2mIEuytHX+qm
9VMDgO8cTSVNSu5Hgi/spExeM/lL+v6Bd1bxPYmrlN245W8jDixKO2FSym2BB1vBuhCYrN5cihb0
xw6BMJxDVkQCRu6CaW/EG3V4ExJxRIZIzI0X+WnOgDHICEsLsUlu8kcSuabOEfoVzXqahRUaTyq5
JPDFua9SUSCrAXRZmpuxTxMMfWPF3cznDm3vwYKNPD5w4Ix+CqogNQfmsCIm0ChqC1uQ3eFi/o3C
U/GHvlE9n5JijmgyDNFss8+l/KRZvlpqqFLJMIi0vnxroRgkWaWPjZmQB5GAV3B9wnyzbdJB/N9B
NHNhwpusEsdlAdaEcDqqYWq14h3wuK3JIjlR+eUwHR9oX22V3OODHDAgDH5KxAqLG/d9cDlE4UfO
8Q9DsPJ5U5AkNUJhVu1ZGIbnCeFPKelOrbPzS5e05Owfk8L4Fm/NYQnCa3UWgqfupVLrboDfKt9o
kYkdLCnbqI3B8OOL4F+AozMaa4/lWPXMh53NI1LQee0AGqKrS2kehaWM+LwcMVcpXPbGeszC9cYG
5fMmBPAgHgr1E/Y2uZgi1PXNLAuAMQrv2ZZdsP879rAuorM93iWI7kUuMgAUKMcYyyLhpCARLHEQ
8U32QWFr5rE3clGpQeUMuOJs467HUZGKU3kAmI8KE9AVi26RNIvbftJEj0LePZMz+Y3oZyXNurrC
huVGcU/8rUaO/bjBnyOyDg4FrYYN8aTvVbEi0cMRYLyr7sOzjKtJR7NUQFSpM3XuCkJiD3dKgpZi
0krKe8BG75XIMQDhCMPZJM5VkOD09yDN5UhD7+zE7oMCSg8rJvCOtDsfstE6sr3eIpsngO4g0WRw
Y+If43R8/DGMQiE7Uv6culvwq84lRzZSwNUCItdqe+k5cmPYnvNcBJ4+ivjvEVp2lULy+uYGerK9
7nL2YYYtuYkPZUivxmxLMnZZuCPY1Qh+0WoJFyXNoh9kxM8FFMPQqdpmR7OtNmvS7dlxfZCcD+1E
ydgCaF87g/QZ4ZgQtbWCP/SPkAxwS/zpk83UpDCGSNqWNyRZYIsfOxoDJTfZUPDhHm7cQAJpQrjX
smvr2NSSiRjRKdrYDX3oMhdCJLXMPJ34adRYRj7oVfCr95wLfbyaaBL7uHqOxTzncV1Y+1AE8JCs
tjIS4/dw3LkvVBdcZs3CbQMjuYE+5Hg2xEHnvaE6vrqSWOEX2a7w1USsbqUF6JzFkEU9Gh0Zn4pE
OSw9AgbCQtkBkLaAtdQOA4EmL4kQZ72OyYiWh3cNX83lwBrB/iZQI4yhEfFu6fkxup0tro58EfYE
+w4CnJ22YKZ5LSL/DVMjDxlStzKk5yB5N05WR5bvJUHA65NwkkhTHM/4b5Trtes+p9FUlv9dTQRR
AcP4PFilfCoVM+DuDBy6nJWx0CXRYVTtDFbI/jyTfj3quQYfM/bK6+oNqdCBgTbDvVhde9+nBr+n
DZ705WyN4wZ69pemjA+oMQP8glVNGMfetutuyRr0iKIcGOREW9wWUqP1tyiW/AqbOLZ6lhh2WHnD
A1uMkOVsf61p8TuTC0qsjqz0lEGNPXYI8VC1d0sA6T8HpMk3UuA7xH+7O7/1xDDqsaFAoobo1bOe
J+Zs9qlBP7tZkJgWy3QKcrl59JV25NT6Rhmiyx4Np/9d0KvYXWxwVosTKC/DOE38S9T5reNKZiyM
pGOumw6JloFsVElSXuYC1fjkwa0zMXH3Gi9F2xDMj3LogUpROyCKYtAbbG+uWPlmBYOrXo3CfaHP
riAzh6DdSTOGyQKCURntZqaHVT03dIZ9XHHtCQ9B5oxuLhThOoqJUBgxPzPqrI0CJKiPCuZ7FJVO
qRDv7XcD2e/dbnSeE99NyzlKQK/ML3s27oMOl9uEIYHTD27oQIUFw8IuCFV2K454tj5X1lYf4fnA
lTzwK3VrZ1PooAThA294+YsyZFSDwK18IgnGNVvVbocLUphrLmlA3DmPkGeZe1pao5rTw4MEFXHq
g9AyQys97y2m57gqqCEiaoDUpsBZznpyRmQOOO+WhN1ABpm+EQi8lVlore6MA9UNgrlN0tT5S9DA
idM4Ebx8aDeE4BadEyJ1Cq0LXnwVSIPFIJ1lfCf4+P/NbfpZEaDNqDh6ip4bpFXGHHN2iKDqtByR
IA0L4jsfE49PK8nYB+blS3NAOESJUm8Brjf5pLbQh3L8h1VuM5IxRcAUUt71QCoptQH7WDuYNtmq
+KCRKC+BBXQubMLOMmCVq6k0cZwj/y6+opPvJbmBneZEf6M4eeTEYoThtYgImmr2EAQ3WwYDinnX
1eSsX+7WFt8M6E4YO16pd29yT+0pBhytiu5R+Q7WUxaUD4DW+4Mm3CV+7LyF1hEPrEgw+UQZF1F6
t0tUy4S/8eaN5wGo3+Usxku7dkjFLd3Ci/dUZZ7xevAumz69NA0Qu+RnHPVelCtN2tBEa3cME7Ve
wz981fd2Evgxh6kFAc0CogljPKNQBgw6mMB4jV9Wg3gcf54xtau/j74j+AsCTDUlbVywZ7oMnA1y
XIMUk2OQzMWRBebDzsUFZFfLAcPVxxcXO0cfP52e33ji1+yna7GG2sEBXUM+QgDpLhO03luaTCAc
d/igllbeAeJ2E4w1JVfvlTM4Exyo7X9GvW3Hc/dg3H1WX8A4imuKZAMh64Gcs7pbZ9JKmx70XQig
aTt6pbKmlYbRw1h2k/Zp/W6uefuy1ROnbRhNt36BRu6Ezp/wJjpw9+UmtVCyTSe21b3m8HYeaoVJ
01ziAh4x0PDooEqxj2xwrmRxmGBIaBivrUI14Gti+rXBsJ0ZcjH7PLZWtyp81foBNd7DU2EaI+WM
Q9TPQqAu9F5ZOo0tN5QqPdeXJZtizWMRVnle1fKfHgC+1ksCm1BYFq8V3qdVIX6EZOk46s2wkPSl
0SrM+fr/NC2WsHv3/33DvBJ3kPruA9KJscAEJCGHeF7bUEPmXwMbdiPnMySPbjwQ2usQx0NFtZKF
fW5uR0ggbw02QpaZAl1dNk/GbfOExfmZx2hMuAozliWkkDPD0QSiQ004qwhJGiuGxbClyYw2D82g
jX1zT2cU+VKkLFkDmWgZj3SVQAqflQr1mEZTh2fcgyQy0XbIFuEbFqHa2vcIDu9ywMfcsyyTr4Hw
FDyA72JFWM+34bIERewdRak4vQ6Gb9CaFymjszrpkGB2NgIP5QutW5GdST6BJbfS/pTuGrBWBwdn
agaag5hTKASxh7QqDuhZFgcpgJf4NUhS6GafNbOTkHTGVO0newYm9adhV1ZPov+U4gSjX6kz1EwT
6SBH9bd924BwpN8Z/4+zbymvfA9sKd5xo11ebKTF3SKR4sPqIGxuYCTYzqL0A3bOhrQifGdwTG7M
9RwoKwvUL/mQxHAByJ+Zpgp1OFEE6pggf5voJlYCqOqb7D4QpamlKjXsxY4XKMTv0p/mb2r7gcL4
Pqws7gxP8MMK9jDHh1NwdDyV71Xq+E5er5uDtlRm1rUEt01fkZmFlb6KG5kcn7nmS4YgTUASM3pr
wlsLH+FrGzHtfNjfZ0atlcbivjfUBhKi6mWX3Fr2t7AbhMYIFe1UY2KWEPls5WScpcCG1IdbiCf7
TUaQY7Fb+zR4e8TZ5p21NDLPaVyANt6/ykJDJ6tirECSEiIbJiMpCRv1RooU1S3OuP8C8qeJ577a
a2pwPc6mPyY2aGh1jChX2PCFxIGWuPPMQ+PJCvJFx0T4sGQFcyGapMeDNHJyM/KkE8ks1lEMptDZ
mqMRpfDKjxJ/fPNG0GgroYzwqEZ37l04tp6Xnwx48XpfrtFyNWV7HP9xctxKBINBRA5rOtV3xCzj
wO12/57vSAPiqKDFQEZ861iZH1v6VBG9KJSiTAaJDuxYe71YL/B5iNcRCcak0mQxUhvAq2yQ7BPl
i2XFTPn49ySj3Wlq6Et6LF2s3PdPzrOJvK8NzK54s0i/HNfeodPsd7c2BBQNT+nXpPb04L/WacUG
9MxyorX99yqU7r7n19yPnpktIYQu26/97YnSxXzbAdJxYaaVYrXH3FqX2PY8oII4ju28kjOcFYeB
CCZx566nCdKO/owdW1uSyqQPjCygPHnyvrZGyT18FMsDv8jmTeR+R4+xlRGcXEhXl9Y4PtElogX8
aD8WWIlccr9xdpUjAeRWzajAMzrx197pqD3r7aZeQUHsTr1eTn7jDnzbFUnqjJsOZQA+P+xAfp4C
FbBLzlyDoZ/OdcijmGVXl8WSkMVbEwUigeTlpUVb1SmDfoFlC+FKYSgH5c4ACc/arFdTr7PUis6Z
LZQHeJPsg41ww5nlX/K6Y19+IBdIb32eOV9ORYJpuuvnRNQrnFSUdOgdEGTslY6Yv5bRNpzZJXyq
gm4E0BuVQg3am6qnWRAedfU6vIVll+t2qT5zm+hdPsPHJzsH8QD1t2IsyZOLwI7Srw/7gV77wYoZ
O+wg0Hvt0OW7UeaIkG0jwQyFiOGgqTNEO8+iweyo1NrbtatIPpEOTaTRXhii6BSMXvNYgSVP6Ix2
hY1ixD5rS+aa5FQ9DW0cpspXQ5vUjSdWGKrNWxFgmrgDMJQa4VPwyBi4psvpu2SrrxWCKzORVyIb
efIFCdOXygeh83sgGNeMoSUjwVteNN4nmy5h5h9yJWMHsiA0rAON6RfnzOGZRapobcIOC6iOMymr
KvltDW1VQXZd+EnhiDG1tZhJNeA2ZnTEyotko9RY76sZt/8vFw+ZvoKeSI1Jq4RzvlV/s75lt9Fu
sRcILlS6LSt1AcLEDjBj2jofWb956i7EYY6bN0vkkIu9f8+Sbh1sGrvibCHEMFjHy8fkCbaeJuCV
mp4oANGxPUR3hyGC8bEyuHjaehLva+MHAnJk+OhT53cJcxEEbgdOtetM3F5y9ShdHiHv2CU9uyw4
E+nKC3DgFhrFu4YOhcR2/j5Zs0ESkGFH79BBGOI2qDqJtRx9s3R0dK0bwW9W6LIeDbPU6BRNQQB+
fiwYJdvUBwkylBod2zoYxNLgVyTf1RV2GEcgMj/W9FdQI6TC3ETWl56l0n4okOy06T+wv0LdC9nR
tZMYAjvuREQLAjr/CH3ht7Zm1iZYHqB6rMaisWYlLmwHjxyNRXFgGmBNS9oC9cLzzm1eqAGqG9RO
wzqMM3OUkBPI/v2cLKybb/06piZio9ve6GaP3B1VuQiTOR/Uf19k9fdRAaJcZxX3J7OeY05wz64T
dW+IszwaIwpAW4tN5/8/GFPbYPzRXCoWiQ7EQIbBCjxePKKFThi+eSV50Nul6jqhpn1NPqGH4ifN
dW8A3L55x6VX/8B9LCoezA2d7Rl3l7PNOZPR0X+xWMsk9MxztJLx4ssNW6Horu2NsB7cfrcpNFBG
OtiM23spg8bJyeKpnhCYsWHQShkhISIFozkjHSYBIgOPhKznUuO5udJ84OPMC67oSao3/DE97YB9
TuBS5XH/RhMOaigQoUz7R5cgt0ZFoNdtF5oALiRXmcmN37EQs0TAtfxRY0Bfhre0GwrHKogJ2DdA
Z1I/vQm0EV+q7MMImmxfTJunMusFP+YLiPzUryxklT7ZEcKxov0lqBKGCazDzDnAj8JFs0mqqxv3
i35E6uRdCu0aqdu0C2pEdMl7H41yt2ihZfJ4PUxGLSt/A+ytLaUJTx18dX5AeRPbFwNzBlHvwuOm
VKMNhRiuzZBdgNKh/luhfw/APfD/msT/RtrzKQ/vFsw4Nzs7YLVzHz/5ryy+8U1zFHJHHE/CB2tC
hhSVfE5Rq2F2rFgyUuIKLdtwGEQGUJU43CDnsPLGOOfowXqZT09bmch46HXRY0QWRuYUmkVGu7Xy
eDp+fydBLKVtGfAv8Fg56Y9xRUUxi1AkCh/EhtWWh1fiNFeFagihYybMRd4IkTQDH+YRurPu2FKB
zdirf2zBtWd8Aw/c6GEbMRWVfoIR2OV5JAvr8s/txzr2gQ+WPlMiWI6Xlca1KPVwc6v7AX/rGKs7
p+eNuFtLV4B6CiThFSq4As61NXw4RQIRAbZC36jM7z61rubaL+ag09uFgXxEdJ0FOsVUMlF1ThEd
QsfFT8fSLl15WHiB2w7aejUhDYK5x21eyBiO8owGi6+BVt52kDfaueXONhbCNIMQT1+1tpWOW/r7
PgmN7//Q5Lh9yy79zIEdnACMJ0G/KdaK3pwSnBgkm9q5BNFDpnQ3Pb+Yzwpdd56ZEvGLKAS+/v7R
G6tOfR9FL1S3oVRv4YqLcaHPcEbPTckg/8wMMX5ovUag0z7XhISsCjz8PURAHw/Fimlq9mLw5MWk
QF/LOaOap/G4Hu8YGd3OUudui/ogXpkeS6ad3lNZ3hWksXnAgU0ETk4QzBnEsMhPk9Taj03H3FoZ
qUO+zJYNjJNNAedyqDY58iPrJ7tTqW/lR6OUi9Rw4gH6N2LyQglxVjNV/JZkHJGjb4EKTpvyldQC
S1E3mVodQaz3UK/MVEmqQlTWfRNg8gFnP2xw7p7zRkaBljWgExPA7c5ZiapTj6sl+6LAj51Ujie7
DQ2sSO1/tUZOrnsCuUHxmhPDtxj58tgLCMS7I5J1EvsqXo6k7knrQ0+XQsn0WScN5aJRhRSxOhh4
a8CSQ6bEyHKu7aRtOqI2dv4Te8SyvaeEDAzVv8x/VUAigWU8Gwc3JJj96tZHbn5susJvcYKW+LO5
YqMoiRnmvl9Nku2a/a46VDqYX5De9iTgpJEc9xEI164gYhPpr9G46h6mqrJgY6YAbu4pr0i5uvLG
L+R+y49Oh8cGRNGiYn/PVUnUVtSburHweBYmzZnNFlAixcGAENtGRc/lTamwTIPl9mk3XUMA09Yl
NDEfxG0wJFZp2VrnGGDDgIsZE1s9DRu1LxOwo9+lVxYEnmYIUbC4DESz8pj/opM+ZB3NptrQqXVB
j1nZgTXWo6kN9Q2L3ynKXIVHcURerY7MUlSV9ITD7g9TvSuxmSVKtD9E1XX/TQqj0CyqNLPh1Tyr
bo1AAbv5zo8JsQAfT5s05R8zqIEdsI8R+j4KV7drfkKPtPafu3FnALGcw/lBdl5mp+2dV22N1apb
6TNRI6HDj5W1SWyNLH1zfbg/pGIdPGVxvZJT8ncrJeVdic6zDPtMnxZXVQaaMUGjudru1661To8v
Tl2AETqnMDYq66CulSoNzsOfoxLGvZsIU8n3diOqGTh3ei1cuwODSS6Xtpe2cRqHa6kZx7qhlZ08
wvX5aXFzO4+4UswVwVZc5IbnevodY9yuEy0U5SOojUc6wMilHA3e6Pu/dHz84Qh6CUxTgr2RPafo
Zr+/o90BBz/RW5/0cazMFDWTiULTzTapRVtvx6zbdMpY8rbWnFTwg716cvHkeLfaMVEWZfH5S++R
wehvMK2r5UGfYGesntVcmfQ3FpJWgOwZkY2e/1mwWXyNyGuagRLoWE9CrMywBP0utvNWqCVbHvKn
id57BD/wmpyy++qCbL4WKopxIJezitEXZQPDz34ZgzpE25y0CmP3TUapR/+uOQhfd5lu2tKwPefb
G30liUxEdxXh6OjTzemRLVfIlInbQzaWgoXzDNsuu7GWZ89B6ptr8J+z6kpQNFGokjpV0JA+h9Bt
VcDubl6FoY39ATzsAtRsJIMzV9Aj05uPF543805RXaj8pm6awb0X7EIEOIgXlbxVI/3EH4QQ4skO
3KzsFD/1kjxb/02BhZRa40YSSlgD7ZUR8knpF1wxF8tJMF8yX+gYofuWC4615lJKbBUW7J/R6stz
R2/f42hldLSjdtpS/82+/lE3W50qbytMz4Uq8mzU3/DCNwawb0mXWCQlm72XLEZlFXQIWSDZ8hxo
d0Tu6HWOWH8LQtiD2r9mUZl+EmPtA7SWngsy/0DuBbA5hSjsOeWAyhGzMRZfWqinYEIVFWewiZNL
hXFUTouGDU9JeHkQunCuhF7roUdS/hijFyVOWlIAp+sZTCoOVKSC5SmQtQQZmLbj5E7D3HZOs4Yy
487YKq37L3qkogbkpGFT/vL86n4Um+fWLzrvj533v++1GLvHjEGq1EX7R2ZyilT18WjuSQAyjlxI
xxKD4M0SiEl+10WqvG4NImBMfxIXPTnGoLp70VD5QSKmRIzB1EVs32Iv25a9rBiPGGK0TMzr0SRs
IpUVs/fq5dAExwsRp42lbWy/08m7goe1qGFwtbW3dw6El8ILC60P46AhAt5yPzs5U8iH9HeAt/g4
SpRegHm5JFgOKhu4Ze1+ckhdgWMie1C9vyPUIbnDUtGaI2fdRbW/CdiwBYGEECkQehu/Vhx927Zp
bY9v3ynJ/xxhXG4lM60Mib9FWM/O28hzkSL8VnSNPN2WIkNKTT7QuG/1uh+mBWVsA/RlLR6LpRJH
VuYRV6HjD/Afyxreh13ftQ10OvqCh4lEaX93zjEPVLQ0Oce2V8/1v8xCWLxDkyq9evG1HEXhbyay
/WJo9rhYAATeCKbwzoA8mtkkPLt54rMcypBtLUeG9dskUql3951tAyImUzlFo3Z37CarPhyTO0Pj
XjDdBtLD8cMDyUNdhFHqZEF40lL5M3cMExGV4Aftnpj8elk6P/MQ5Y4FDSq4gE/Yby4vEuDPhZy5
H/zLZILgCvJ1CsNJYwfZXjuUOusPhHLo3LDOa0psbck7GVBhbDkcYbAEy39v40CVls3y9feM6O77
+lIkyj6vZSk8B6SDLTFZT5UhyUNxevu3pSshLh+d4uplS2DQNMMZniW5BiboT30ZI3xmUQjF2XiN
M9myM8cGF1I0U/qJclhkkKNhDuDxOSh2p9DS8+hFW7N5sBrjnMePe2Lfn+yH+0whbKKzdBg5+hwz
qA3fBo2z4tm17wnU08NRqTmwFc+SUFw90rkhvQPPsZ+Pq2FqX7xNFDjTG1AAPy3bHVC6X8lW7OvF
A/Xsw+S6VZJG58NY6tFdqYuBE8p2uBTpVKcNSSvBohhibDoaocB1bUplGio5p3evSGGpbscDPgTu
sneMNK7OtvVKeFS0a82qsfnHY2iu/DyTmL5eGOPBACv1NBwGSRpntBkjABQX00VKa6hFosMhdhqY
gMmhtjJ9c1kc76c6CPCrFYOqitDkwkLN96k0bGQAt7sQNSVJCsJIXQvR/kz8LrOQZakx1F6WQxQA
ACRuvOADdroaduwjQ01IWF2ZlsNILOcsiy53wdqjRfWV/023ScE9PoR+lwdJfiZuDoOLXMCKiGSc
IErdEyQvHKWkxUqqowuY9o/sGvJtMmK57pqvhju2ZQUMDtADMFXz5AHi8CXMR/d2l1ymDyAsdGc/
R1e6N3Vxr6fbyn/6cGOBBa2DHnyP0iWOPFmqJuk3DlqWRsnEwaTn/7TqwH4GqcgKIlinVxXJO19Z
6eC78N1O3pYvaRN2xsb6gaGIx/2qcycQbk8k1Q8Yk1JKewNNTvo9X1AK7mNHLqgViw0y5fZdLXLo
ZbEbyQzSnwlEUTGbfmEPdYh/99Gy1bcoNqZypHsViDruQlZwjNFrS3Ila0tvBPP2APa6QU1nzmJl
i7VuS95407E7KnidzTR2k8VhQL5FhCB52a/XZfVCs19FXHjnmPJ7aRm1DH7O/NKDAfJLZxyKTdN1
9+J/IkjHYzGjqnQ7W9yUSC1J/OhMmHbTzoA7owwJtwySz6dEuppYeYzF6FqL2BvJ4JiO2uakuc0z
ox/l6kLJnchP+mMQBXdLcV93sf61XJo9v5EvKKUH5Y6H8afzOZcmCjEKmkFLAfTpMst8UbyIcKC9
J6AWsOpJ2ez3ZefNS/R7qc0OGNOSbPZ/xcdmFZ4OwfWLSY8nNbj+ECAl7nmAZLxE6+jZ5F7yvB87
bg+cjHJKN8ZXz01eZbaBlqK+Ew/V2b6xjBHFwMOTwNtYN8mhglEMORu+sTRD8UwH+lLcDA3+iG19
uFsFgOi/f0TwmxmZNcA5ej0VvKhLS1I0ZmL6P8bGZ6zQKQhmdt5z/46PlUOMV1bR1u7FXuC5kJHQ
KYQMxWO9tCRuyUW6DXNXCVA61mAFWkgro2TvqUZ+k1pR2n5Tw14x1wY47l8Ali2frCxpjaLqpy8f
A7F8haFAhUMeFb6X5VHVfeFguxx7zQ+N4hjuhq3ec3HPIqktIZmMVM7wX5cpZ+khHiTaGPiaY9lp
+6AYWtl1Cvmaptqz5rbXwn//OfTOZ9R3oFrbYXVJbg+bhS3bKu2ef1LgjCby5iLjWyLU8wHOChz+
kIANXT6Ir6/8iL4bw5EwGzy0yzO4sxN5UZmLCSQLIUydlpDrHNiOHem/q3yL/lFB5mT4e3wF7fea
AADbQkmPOcDcPjivABTXQAB+Ztk+gAhe8Gslv/9SJjbRH6u44HTStycbGiQicDk33eTi+6GN191V
XPl/RyNRMMLY3qb/zNKH4x0M6kvW3fl7FWpr+00Za1hcdYknJnHsR/7BsGAuR/OCzxapOp23hvIA
wR1gmNsiMdsjPgeJq9kyolG3Ap/7QyH6Fq1inmYCeIjztgjFqYvBVtL27JLi+FgBMMuOwIh3DjMg
QFtkGYYUfXax5uOKO55d0bDCyA0OcHuKQYxSqIIOxCi3NmVlthHLt0YURn/SnOFRfIvFPRV+5HzN
S1K+uS+W+Uuf7TplKaDbjsQ+LLgIAih17klatqNouYkrjExaxJVj6j337pRRs0HJcZvjhVwhE7IT
d9o7r0ILQwWsirmi9pxElXhXYbSga4YAZd0Pyql4TCKJkWZPHR1qDxR2B7SCZLowF7nmK1eYRRVk
QXkq3E1GUW922GyVmVBXIt8+n8MhkDEDEGscFGHDCYEbXjdxeASfPWAFkwZsJwL6uHFuELEJ10iR
96wTHHSl1P2pxy7zHYLLM6C1L0x3QQ5LpDM9ZGYTyNGGXswDpln7oa9Ethr1XdH6UZJLgY30CNF5
g4EvC0Vysyc3bbsJteg78jxA8aaCm5oVOfdA6mpnIaBwRQApZcL51M9YqVptJyuMsUSaspL32sCO
9aV63YeoKAR+uv1wU8WWUIxA49pRBs/QwlMqcGRfHiNBNQT3256norCK1iD9FWeFLHl18UnE+K9A
Za8ShtkVYjjVOU3mWNbiZ7FiXOXN1imlPDEgNBotvW3OQyCBBnsKvmuBTt+Y12PDMCIsC++2Jp4+
dcqFYK3JGr7uDjBKz9QfmrPiRA2TtdJIKn/tT5ivukYKldmUGVK1cGNYfEAct+bm6E2mua/+3IVP
lhWcu4sW18hBg2UKiEf6WWnrR6qQA4aRggEeca2tUMr3balD+qO1QRP4v9rpG8nC7RrrkiDJPOdU
Qp4VUnvEn1kr+u5ObaPkal9OhCU2T0iPGzKjuQAcWKhymM88GH4s6zg8GUytOlZhxVmEsDL54oTA
9tqmQZM3XQ+jHt7tJVkvBHeMtBAzYS7BL5Gh7ARUcr9Od6BY3vbweVdHLKYyeb5ImXUWxhs7P2Nw
er9SLtk3+kga52BKPHoBcm/qSdWXwOOh2d6I+4x4NmRcK6eMI3BZK1eAAi/JxPux3oZ/TWZPoMKg
JKK3b8l481173D7QHwUqhmbGNVohq6oFaQq0hf0/ynGjLAoucGEVUXdDe4TmjDTBBSYeMIoY12lN
NbMKWDObGN9Dp6F19ZHOOmB5tdmWf5flbCV49bMhX+ZFFUQ5TKf9EbXSUm1o2gBxOTj+2ykZcdD/
Airn6PmD9kwQIwe2lvKwpK2Rhlaq5+jNsSpUcANg7nks70kmk5G1yVbhQ65h5nCXICHsU4URftP/
/1X/1DrWIii/6dCmZUVPOZkruwodZ6bXZ+arzy2UkU7RYX/XqSnertlkIgZ0yppBGladh+vEdvo5
KdCMIX7LP86eyePNemgZR96uAWHDYxDMytdnarJO1VmZ4hsIYWwj+t9+Y39XeGErhOv5n1Kkj92J
0TRnVBPbbuq01+3ofZ9RNikD1G0wAbwT41SxN2JyAfr69l9u30ydBOXRCXx1RC2QydwGah0MLot+
1GYdsZ6jtzTyWIxxSK6LiasvkoRRFj6BArZxl7ufy27Sb+dp102ku/v0j4zgiVhksMXadphv+Vkj
n+0wWnD6wNGMTarf+SSfZx/l0z7nVNNvf4Eg7jjkhMVfASuOZxnVHZKaLcm5uqCUAMKbeNi8p5rE
GfHfM7LfosdAJ70x8SD7phQLZaZd7BISNBX/Mc/bLrvzTQ+ZGq2xNnPEd8yhtush66u/k7d5Ua7r
o01n68/hRnte4DZtRigUHgxibqemB7WroCeDNPII1sJojMVDo9C16JHtcrK3FXl5V9SzAx2mUhox
QTaurx1y/dGJCVdza3SCPclZgBJmiU+DgE5PkVKcWNfpMyTDpLyqmRycmf514GGAjZjxpmFKcWiq
TTHcsUpZJma/bmn9AhjQj3TyTNM/UV9FjXfidiSvfMiHsvm03EFJYfShUsDK3rSSLYJLsHgCyANz
3Npon30UyrRD3cOLxDX32KWfWC2SOHGjwAjRkYKwhcSsTXujV5HOixlOkXaOe+Lekis07N6tJZF9
n2qWR8Vi/Hnquie6BCeHRIm5/biX8SOxY/gFyla9BTnnyCzRAoP55MQJiKPJ/Y9uea+E5Wbhy4oe
Z6nLQin+5QYzjc58bHTrswryeB135Nx4A2RLq5khbNOuz2+17hmQ5QNOTUUu+ejP8ZYvw6hpBYf6
KSLTxH8PdiUTnhG4AUSAqHDCdCuV0D6523QqoqjI8x46oO0GhaeFscLAezBEGtUBW3Ib9yW8gjhS
FyQd527NM3lev4I7HPwV8C6faW2MA737mmi6lBjXXIYRFw2o1hvVeZtbQhHqY8P7PjfGTV2MToM0
D82bn9RPpstNLZ9sg3HFn9GOYQi9ccQX/L5JDOk1u13aDSqMEoiT1l4BxCiereESEzeiBNB8R0eB
MGD9u/Ef7foP5DKqwVKuJL7yb9Mn+Pr3fTwIlbeJ3iAdgtZ1wZ4hj7q6a62rk17shJLZB5Gr5YsJ
R/3/liNU+L6d3ap0UGp1G9rzjMpploFEYVbJ03ZPtwwavW60Kb2hMeclnZ7hlgExfHTFtFqOMZ3d
vs7FIWDe/lz84AcBxiEy2beYow1+OhDPFTRgq/u0FSrP1kwN4ztvqFyKtoubYRg66w7saSc0qr2B
y+186nGcVe71SRZFcUh0Yl+T/x9oWApGyMKxicEfQs4KRoVWABEM61OH48FLiTpFfACegc7cgcQ/
jG0g6AzOwsrpOlgaH0Z+amyf6ayQaMjL9I72gpDKZCHY2JpymaZS0xk3faLNYHvMcrwPfcF44g4s
bUfcBb2G62UwJUoJ3oNgfu+EdM7bWBXJPGH/SpdOUq4t7bIyXwMnjYqL6+Y+8pMDntN5Zxvo5cIO
X/vBXEmcN0hQRoZNBGIigIK8hjYA0trqdSoJghOEX0TKeCACz9FopD5xbD+vongnFsSdacYJdXbf
7DO3C1bEn+L1GZ1firY8kJzuS4oXLiZGEDE831XLRdlScV2tkbTRwYSLXIf7w8/zV+4rJAA2sD5g
37hvkSuPYQTUw4AKASj1RGUrinGa3H6tT14SXk23TPQxAbh9+n5kvu0jeeDTns/VIuF77nYhOssJ
00jaV7COoLD9JWjGBNYWVl4n0LjUTXz1POaFe57IfQUV70Qbi4k2F2zSOv/UkL/Tms7I4O+b1yu2
pH0caGAXsTc0qlAVq1RG+FX6SR+9l3sgbGrTPPoIw1tyzOxwdHRtPkH14n6KWdF0t7Z11oijr0Oa
JX58BKhNCxWE/ovqi8aeYsdMlnWVqr87TnE5pn4oOKhbb9iOOHysIoe2u9KRswrKNFFb4hCaP3n1
Asp4wvhU+qKt9NIO2MiftIuIU0VAR/ecsDKinLHrcyMy7M6qBdfSRDtxdOiqa7GpdSpVDtROcw33
YRDcEvV/lKpd9OCt2putiO8ENnTthyTeeiJh0qhfXQ/B3osIo4oPDgNBbVRDJh/6Nv+tj29OA9jf
2osE93+PMji2HRpCs2EYytVTeqx7njUnMhTZhOVXHDFaFfUwILdP6BPQpSq3GmncZZM71kjVCPGI
l1x/6MR6k16ybqbafZGDGeQ2u9N2MhcYd9ChjRm2HMFpRe5IxhxVWeKYiIIdAT6GrAyji7t71ub0
hMDTD99zi2pnAzxWtuOsme/04yBvOGFGKEwdmi5Q4b5XLZTshmUaJS+kNhfhQG7KVQ9PoecE48G8
gxfj8ACfw10HToy1m0NvG7947tK62v3RHVXw8u0WcM8HlgwAB2A+UQpNGC6n/BNLjxneJU37oOyu
NkB1F/RHdCf2krTb322zcIFMYk66rai5vDOgEB1DrlPTka8iCYwvD+AMUobOUbWWmPLnKw04xhNc
iopTfUDkMr35f5aHyjSHl4i0TSQ3aD5gYOwIqcvWjUHr6QLB6ijBMSB3hDrzRkwa19mqTbv+Y7O+
ag84hiXd1+B4cqwBD0XZJXEi5879eYUDa8RgmoWMyWR3Sj8dJHnFrch28iUA01s6lblXwD9kxoE2
Jisf9jW97DqAxiSsi798Tk9LhmToTQOTpJeJ020zAoff8hc1E0wvL1XrBwQLe5boIVoRI2Z3YJrM
VXklKsQWwxjJSSH6jTwdJsoH7M6qhw/UyxCWyZQsWA4Ad+TEcmmROsLfUWdr4YxzIyx/ZMUy7oSH
VXctg9NyJP7k+DGqveRULxv6YKs0YEuceWRXvUInOsYZj4my7jnyNyKypDFi7ULRzAU/t0Qn7uXm
Y100EeW7nE8fo6HhB2U1CjPj69M2cezdeT6sPgD/0pvNxxXAElVGVwscArR1am6bPlEfllPR5Hse
2Bwc/VAtWWbOtXmzNtF3vuc8anCndTZjtbLyk8Q5i7PaV2Vsf4AqObwujnWXyofyYD6zQH2wN/Z4
U1d0xet+smEf/TXi5sfuoZfvrQWoH+HvE2aPBtl2vmDCBaJ/4AjiDdvLW6/MufaPUV4ZqkJCtzWw
gLbCrXvi5A2uruN1XnW9Xwss+zx5dUNYZHusf/60ALFOGHXyOIK046CCvTvhvsJPlDD4Uimj2SCM
Bs1Cz2tk1frT674FM85p6la/7/7SCCsx0wv8Wh4M6Xy1XN83lDJr+DSIdHkKGjuE67Vd1KZK1X4n
9QhYPeUn201yAhoplpdEAoWFhzixG4AgHDL9Q714Zq7muHSjlcawqcFl5PwS0aTcCc8orPS9DHaR
ysoic79SExzqQNW1j2Qu2bXHAc9LlG5NwTqL0W8GZHGpD1ULNiud1Ic8M+4hrvnHef9vueq/tuz2
j5jH22n/06Lm+zUI8zgiDHS3lKCp/JnSDrTbHTYRbbSoBohAQFPbKgevBz30RborYIwmydAHQ/nw
6/G9730VgPoDfk2RSUtMQbKGVApa9VngGZBWHadBg4qf98SP83GJAviHN8gR/gM59N439yq+7S2h
tRxEO5xmqkTz/ld0cPk6J9GHdg0hKtd91l4P55seOJ6+x1v7FSrkedVu9LLMVmh5ffuEmKI8/BoC
C9QHjtEYEgvuKQuVrDKCJeaLGf8aBvr30qxkpc+/OXFiFjybix8joeyguyC1HUpeGhof6zjBuhqH
Smr5gUjs6cTBf9cK0bXL7wz7/LoBc8bhLZ/bmXE+t8Qlqb23anUpgb0n572P/Ued40tyuIfCbaJi
/YcXdHhHysln/9UFOVnowJKMluyy/By8FGGpMQ/z6u7Z3okLUqUhzo5ZkPqzhFGfIwSg+iTWVekn
IsgRGNwitssaCZnR9dHnse2ZJLcQjQfFNZ8tj1aVuaziD/jhxbCuq7JMIdyJuqK3xqSBrwiyrJR7
m+1SHwyualE7Y5/BZ8kGqdLqy4h51650PLe3VeN79U0PgyN25S+WnLiFkjAfj9QxyNEjhRCkOrri
pqTWD8RqfgAzeRh/cTc218XgfJktjgPH6te7ZYnSpKWRs4B/oz7Wt4WJnykmv5a97XvdfLoqYiLr
5Zm8l4+Z15vy7luDMKZdqS1gkUtE+A/U4tgupnEpR5fL2FK+EPlMb2U1Na60O4JQoTaAc19yNN75
TfBElM7GSf09iGt0Eq0EMjNEBjGnf2gNFsHol7paJNQXZpsZ6oTtIJmsunz04LB6he7AE3lhrM0z
g3SONGPxSAIDw7FT4zCb/Hz9JYBCoUw5j3YD+wvcMnQNIGnkgJtjpoaJ2VJ0EMpwmKs+K+DEJ+QI
mc41hvB6LGQGTwEKelT3wTX3BhvAOwKvBb87m41NnW8OyA3bCe3TgNwZPj1xVnyRKchVV7wFm/MD
tZtumzWJ+zFoaNkBa5aCRjRBmZrCPR75IuRNMUqRHq73j1X+oAC2KHXSeL6CoXqZ4F+HTI5VSx4b
tx9ATaSvNrNPp3p/t6XGi+71MhO4iGw66LInN9d5wxl1txA475Z/63nJK1VE/yuA2nbSh1yyTsEE
E1dEgFxocin4srpr1saDOeh9XjRMf+1Jw2Mx138fWsS9jFB3XUJlekzXRPUTpFJqdZeRHvjQ5hPf
Sj+pFkZsthkBPOHLUV2oOo7IZKWbXUrvbceoKLKuDv03Dhhf1L3yNh30r6QwTcz4HDmo8LM5cDZx
Tq8mkDZAvp3hS9tCGXOjKPDYE9wCqV5K/mHQPkpCX3gRtBB+Kh7jGrHYeBlrXYpQHpS/haRvVCj5
Ur1ycz8cD7Q+wKWvq6fJiNuJ/Fj0ZJxi7wrAAzAFRz+/RIhwJi+r7remocE9miZNKc9+DZnCSCS6
3k+jigHGT9U2e2Ifv4dbWs5nVYYpsneWxBzN/t4Y4Yx8wPt70eNHcyjzauR+tzeMw/6Z1CVvS58j
JO9QwXIKp5BnF1vIzmPa4W2rxVieCHBoOhDlvM7df9E2OhJxM+QVjaLjhOJHPlqYqvgBUjRmaOwI
eIK2hHzFfvT29C+1o4yt4HIWJn8QcZJA3nqi+s+f2emdEFLw2rvCbQTAp1Z21GnhEWb7wUu4/IaU
HmyUogh65QpnCiS6Z67PyZ85HPK1McQEHkfli3RX/V6OPAXnhNtNnrXlB1tPfsVhET+3ouJdvx6l
sfNcFGwZdoGPtTIROxUiQoi3Vl1Ofp8GhBzauiN9Si7pOQyQzAdcg/JrMebz3MS13dtDC34YwPGU
miMtV6mJT+GOCBUkksiAzASvo/gBiOx9dzxEi7owtS0zGcBC5h0pLHwDrXAeahRqogu+H/lmEG3g
jqkEU+T+XLvSuNv1CIyVwqk8w9LkMFt042pmvtaNmT/B6pZx2FiOSAynlhO7CpVL4zDqgpMB/hJG
o9GR1MXReQ5Sp2DZhhuX8b8OnqTqmBRpcbdDjo5Win3CEKfDskSdKyXYLkuXB7kQmwP3BiPDD4s+
4DQv2x7+WIc2sYr744hDXmWhKEGkdSusWKIO8w6+d3lVaH6pIicuT89qLpMz2J3kgPm6VhyueeRG
pCUL2Y2Fb0+zq47h1a8AN5wYabAblkyREBDhV0xZH6Mtnhua0iixEhueqETNX1bYwQkYZvkBeX68
1lcjb27/cgMsXZIICsdtZAxaNS+xc2Y9nLZmqiife4G6+8etRbOiYt2GnQUyAIA2V+oDjaIl6IqF
dnLhzMdg39S7zhAOWP1qSCjYFTht4bKSAlmrJE/PyfnQcEtw6RQ481G14NlZ3mIptaOVxzXKGypG
3Ul2ayyA3iOPLtKtoyErKjkurcVarz9c/bBS9fzgfIima0OUQv/RZ86XaeB01G56Xu4l/gurhkXa
5ypwqDi35u/ovFywnumJKC8riutgDhitVSGWr8iK5gE+ZVM37BhPbDd2CIOuP71RQI97kZLs5nfN
wjpA23mFAmre7xTK2N3MZDsz4oACaqpAtilHdpeEs/JYJcI8p9nVZTUaQHK5w6H5RE+JKcC6JsNa
icXKWfMkyRlPY1bwKQc9IpM6DPfTkKRiESzuOszUETOXE1Kn/YdS0AEMNzykkp6cB+tTuX221hdL
5PqLzlInpYNV0XvO6JQ7/HrIoElJ9UTc8pXpvFceMTDM/M196sWNzO9O2YMLF4GgecgKgWJdtBij
XLDTFZttto+uphI9iCG9Jysth/1uiEb9h3eyzPlKs8wd07yVQNEd/aZdr6i582AXlWu4QcYmA0IM
nWWDsDfMw1H69a1n1bXzdcYs7R+ny7UXdkphf5OsH+ZUTj7kZWX4SDRoJfiAJmG/ZFAwLEtHyn+K
f/5B/585pRa2R4AO1SUc7cE8hG8i8G3bF7mwPU/XygL04e6EAaPaYCjvn9WlhQtv8YU5M4/ngY5m
9f5/GVwlyHLWD/u4FU3SpUutkkjUSKYJ05Awd4KKNG2MQNCsfUAL+Mq+cvzSzPpUTjxkyvF2EuBB
L1uwbaskEGbI8A6eEG99KR3zVCbxm05u4ASRdjdEBUK4ve/dgA7CafHtSGEc7QHyYes38/eD1SEQ
B7jOOi9xvSixQvK4VHyxbkxDfRgNGy5s6T/7+kvuK8HfoDEVRI2yXdvC1Jkf52Im94/s84lrr9rp
NRrhyaXlUqry47aNgVeGeCgMoaEjcYiQ/KGTLRAKqO5yY5vzq9Ra1/xlVqMLGQ6LEeDrlIfH+PXW
+kkdAGNeenvZUN95A1DzerlA1AhDY+ubuvXyvwWl0s9CZWk3JWJai0H4WQSlbF6tdI3tCOvCMV12
b7Yj1Od4USpSrB5Nfm3g78mGnOVQAlnu4Vxq66BhWrN87rsgKAPh/P3wItJE9RUTzGvog5/gT9bS
g8ge6Qf2LDWk3+mXR6YrnBHyH9tzUJ9BoCv8D403wkEgEg0j5geQVOrGYNdGypb3kvJIZCzImdsz
ITVahsKRJxHiz3EOirjPZugTW++yRnv1TbpPyeYPgzs+stdb5BorGodS2pk8b8htLWNv4NbZZy3j
7VDJJ7EjVGznuJaLwevBw8Tn2DYD+tRs9NUD83WqsOo6XtnP4h90dc+fZG2jqZTryRefc2WRWT50
PxLkFfIx6sixqYcPFgcUxrNWboYhLjzzEIDVZtIUwEV9wgZRAIA+S43EoEzyHcTj6g0UoC3xS3ZJ
qBLJNbCEYIUPqhezZKuHp0mugrXXdrwMhaIxw7HgvVWM06dRrKMKgxlumfb/Vgnu3iWIl+eFSF0g
FRTFxN2hgIJfWrW6KUJT+3WuOAMaFy0tRXqr76WFQAInqNkuN/CpfSKTCqATX/aywylL+IcYZQZj
AtXOGv36EHVClexEoKTg9rBH+4kFGF2gPPd7QLm2DNOD1UvY2mJYbW0VBoYvRc1Thn3D0BAeIgwW
6ym+FTWfc2jferukAq7LkTuEx1SdA9Mvn16igJ76FEYvceV4rRx872xvOmQM0hLm9IUxeyhFbTGk
R2qG20XcTQqAe8WRzi98HGj5NZwboS+gSBsviBevpQWQuopBeyEcmZbV6y074zvbynvobctukbVD
mRVemBjVEUa9Ml1beVW5v0dTcEk3REMEOuZjx09x83Uppt/Ou2W+dTcufIQ6YqhvLR0VlbVQEw07
qQRvlOwrvyjbMT/Hg0WKcR9PyPz5G9ojWhQOt0+ZXviN920Gqbl+Yy6paycNHnq0UrhXKkx78toB
P+a830orwNi2tIJn8eXidjfEKy4vmoBFk6Mei6LqykJPPo7PSywPzkL6sP2rRrOrgtWN2RzKtVDx
CGJj6zVxIv8ylR671BLO7VaWV0oozT8l4ZFCNyWqTdqoLTeU6irS6vn76K2ivTlbLV1l/9+CXB06
lY1fRTdXqOlywKJwLSFbFZY+7vxUY7ViPWcnbV7KRi4UGFmyjOeb2tn3iqH3WwsRpom4fM/DbN9u
zC45xFC2vrZphI/6uDR4bmqZuxMM05WSsgD3kh80WQ9P/vTZKUSVHAVUwMOssRHGO0EZO4K9Jb6X
IZ7HBtbe+FTriYkW+uRbgszDenginDyKWF/H1cUMD/zRSwfg3feLA+1DP6/AH1vtF19oAhxhEiGU
MqYm02K5RM6yOeaV6QCwk7pGk1/tVur+nWr6bx4sbVZMs/pgm4KHXieQLA0nnrqWAJ4TQKQs0q7f
pl8WaIKMpvBi77ivjYit3L+5I2i5UU2Un4q6/eR+Q+8JDpj/4m2Z9AtM8FBRaZmVfhkngvwT2YFx
ZidsxiuS29cH5YD8JWPYlAz0fhZg/3Qs87SXgwKePTU/OZWXVxANHJtbUThoWW0K+2bMH2rRUUmg
uk29gWXLVt2662ady9FEU2U0i5lYbvTdt5LYqn31UtQBbTnpppBeypVAoA0nwEY/DkC3ejkUrS2m
0qMInZmeqAMo/Frr2Ejk13bnDDsPQbsRq/AKnkh0cwTyOcDIXDIYO9Pa+bjLzJoPU+uC7kULQM/C
ifjD//GJrrxOtET2cHIc+fwmNK6+TwFSUgaANTuApZ6PbtyWelunsc533xypBsDlHfZSOAo/ezvx
uPz2g2OL4dPxsVcgqaskKXA4se6ynhx0eYjb/mVtH0cr1f5aSFJTg4TYZqHSjM5mrVFlwRZpMIQt
hVoBEayXKCBvSPQ1T/+H5XiirqOB73BMgFp3g5LOwoPaFbLZFeGeD53wA/WYXc+i3htpkrIolZi0
1D/U2D92ZrCTZa69DW3WbYERsHf3ZbxlXsStjzpBeSAAQQJPTJFV5uWnKhyyxg1UDe4yAyZo4GXN
tXzK1e082wZdYpkcspYZ98pdRFqqukXCrAsO0nXUkNZzOhhESQXXh27ItlW0srIxhz9gM2MKLfHT
5Gy7oW1wZ2JuX8a1AwwnPowFqSpLiX+MwMuo/2oAJ65QZat75GklR1dJM7IYT+csFRLPxkCVnPbv
xyxWrjj9+lWyOT0U473flrtNfdNMwypMwCx6DZ8Ra8McgvgDkd5zg/DWEHckOfjZzmE7yqNam8rV
0zbWjR7QZwJbtFDalr5SLC9FWIu7vDm3Bl1o1ESe3HOj2qiEGZghT1zJeYBxU319hbUzXulZLaKv
24cL2QNTGsQYnjzCpywZXEQ9Mc770Pe103rWdXtU8aZNH2eTGGzMqnB/vBCmGulhndXLbpv3tQB+
DkdKW4hfk8Rlkp8qaQRVAPnVrRGqzXjhzC6Bx0T9XesVwEB6G0xGleohn/8YyE+nMUVYbSLXXE1P
oWq53PsBplFyvnME52ACCPxZr4pvKRx/qXEyss1REkYwpuxTVQ0KOS9rsejledHZX2416/GZg/8Y
IoT7j6Sd8YEuNtDXxz+TON9Tg2oLTLWf5AKPrrN6/SNO+UDp4HwB+U9SHCJBichD3itbdAbdtS1C
bcPMwT099LTDNxoUwVz47myVApLG/uijo2+hax4Fl9xOy1FRV1DIzC9SMFqruVTzuD7dyLueoxh+
QPn2f7UWgfWzGfOxQ1HfOMJ5IJ819uQKfgXfp0ctQEGwQgdVPKjKiu2C1UHreHx6qn0t0QfCl7d0
tD7FnObvXHFaepzy6eBbkuqaR02+0rM13SaUmpIvVKNQYI72vuUigV5+SeSZI8QEk1Q9es5ERA7P
bVEQedyLfdP8BPUnNOESahbjDee6SYPD0HThqbvMnl+GP2qCgygrqZZcdE0ScnWTSnXhWGQRUtZI
XZuwtdDe2EFuyQYCb+kxNBR32q1gOI9rt0Ut4HxfEp5jUo2RQvsXaNQAAVAX0GloJC3aZvCo8Z5v
JCooVhMQBFGcbKkB5zsxtDqlqtlbZ4M6kLuCxZ7NG2G6LVw3+BOcEZyBK8R1kPhhcjjQ7DXi8giB
dgSIwezOnJFcc7cALsFhpJF2Q/aU2NWfIKNiRL722sbRtFoTPsqVtn1vGwRh5HVat2IDJLRn7Btk
Bp9FyUenTMXLatTkP6Nok9xtbgR9zKHz8WLI7YilnU4NJHjq5q4qOZECj+gbHNN1yd/f/gp5yI2U
QPgH8YNhz8BwWHKofMmH5qxEdrPQugoi8yNCiv2Lp21ryTRNguA4bzzsHJUKRc/Kyl82X5GKWfrl
NkHNm4LdkpV8yLpBtZvmQ59/6p9lAukfQNYC9nsF68QwbJaIYnTAeu/lFN8gY+n6Q0bryA8UGkDi
XTkZxpbinkyum789Fv9CTaD4tmS2dh4d8HyyQ8Gioto+lTatYmuDP8eWJHXMF9RCEu51HZLWMtC1
R41lb0DDBDlBa+fJY7+PiZHgIQn2mwKEniHp7DaBCnampKS0CVsxsln45Wwgi0x+LdsTuh+Xew7p
56RPDl6YnMe1eIG1NVTZfd6+365WdwlT/thXseKBQHCtnSnvYpjK+JJgD6IKBgPSV8OE6n+uHZ4c
p26+l1kvdj15a+vEnLYo9opTS0cDL5KQWHi+QOyeCsI+bmscO81FuxptMZ1AEwvKHqhnJa9lvPwl
abNyLluoRmmH9XS9G4tIz0gegc04TG32HUgSQHi0q9WdCo+lmR7SjbwuFZfulv/T6QPnK4rydfdt
MsPWxEC2tC8GbbM+NefHchNafj/SrehG5V0cMipMLvQciiHsud9QEzAU15thv8Gpkl2O2X9Bkhnm
iwLkfSlll5GYi0G9ciHh5nbtpX7G/lfgT2lBxAhaY/ijIDKMxlb7kESnfjBPuPuZ4L64Gesvd9+V
7fK241GAEMAKlA/Nbb22BazVCtIfPWipYeUwmCL77BmRoCrXC1ET6zAm1YnLREWjXKTXGXvMnRdq
RhVWxx/0jqvd5SyOlTq7bCxSnAmZjRLLeVtzU4MuVTf5eZ11dhenoUzSW5q/ntTnnCrBz/UwIpMW
CplpuR9Tpu/2DEr1vI1CMrFmAeWsHSRu41Mkvv31qFZ9V1vG9QoFlQXPeLAjI61oHcCmezeNtqF6
660ra46WyKSmgX078gQgzNNBYoyS71ztBPlyQChwitg3diWDxIOh3QqCAKkuyielG/Y7NwloNCXU
WKYf+8hyslbClKvjZXhieaSbdKu4vr2sC2ueLeRfHH5lfFs0fvogztcU86MzNOsAUdKV6nlpbyFh
gmMj7KHp9XHqiwPlkAyrerssCze0HVQOGtkIroRXw6G3+w5djR4xIwm0UJeLzZpCXIMsXyYFO4ka
IcHp+/bvXvYTtBN90PkvsO+QKPZhG+GD1xkM6x016SB/h9uHVfMyAamJYb7c1L2AlXOz+mhjX+0G
ZYrUUgnbRuVlVRyj6/hxy/r1gfsrsVxANyxy0csjmo8HwUodS9ZW04tHzHdXl5Aw3r5SJBmPHaK3
W5rnjr9LV6MrITS2jToULuf+vnikUyj3wB9/o2uXU8mALqBUjFSTDpHnLPi2eotFyxGqSvEXpR+S
GMm+YQdwcYohNz7izhSspuhsRfPLVBE52KxAnbSgJ5U+ftwgARqv3BFad1z/Z4WK2DKsF7H4Vafq
Yj5OQrIA/wp3Bs4405gkWsbxpE8yplkbJk1gR7Vpcej3ispXuPJiy33DBaI6gBjafP6VWTgH7FY4
QyFlGcQCbjOgVky4CTEBjxl0ia3pNrwzIbEv0uKWxZIaQwZwMbzi+7/lY1Ud0HHNrx7XC7Rth+jX
tSDKchyM1Q7gRqjcKAm8eQ7WlCX9lXc+cOCNfp5zuSThcyHlgFRcUjBRU8GZ9BeySFZ479ZnfS7J
gCP/8hu8rsZH5vVU5761BArWVi7VxbujNhlznW7DuLc/FtgQbwNgJ2EW5R0WVYqqHTYNfXc4YUz0
2kG3a5oMaJR8eNL/KTjtwTUvxoZPsNirxy4ikwEqldR43dmfdBSmlnvbTHzygHzSgrkKhKHJo1o2
HzHIfrGoM1zfX2VDX/v2vVgNBM+s7akhn4vYCNVxPzdkR8mYVJ8b3HRWEV9y4wqCJjzkW6pYbqUC
+I+xh4Gjtw7h1l9jAFVSLfSWoUZ8INGcM1PHIouae2EjvSyrUr8MpKBVU1lmb9v77HN94s1phkkr
kN0UR4HJWWYFC78DIl2p27wv4NUOKgQ3ida/gVoQgDpTUgeSCFx4aM8zjAq5K2fsfvsz5j7F2TXG
Hgvru1BjpqwOW2i7HxYpbik9cv29eQOCjQwXFy2FQWZX7tV7ZdMalMtyWyiJ7s1hQC747KZPaK0n
QN5MaB6Hh98y89QcUiiXKeVw4gm4Wj0hLA//VkJHdskFpyUK5NQZPJfbkjDu8KcdU7VzpyDrYBdi
XXIKQZxg67J1E7qGWb+52ypQoHJuWLC3BU/cQEgQjSwC3wdr8tsMrlxDVIlPqySxfvNk5FFe4dUN
8nRdHfH5ds3onhQL7XLERX1by4rCff/TcT35VHzTxm8vA8MA/P/9sLhmVQpontwZy54l6JTHAKKf
ObHRYi45twKQ6y67MSHhhyd5q1j7m4t9pfru0Zef/LH1a7Y7zTMaYq5+c6HqyhGw8mEjsPEpxByf
XTWmFcfUjFEwSecqvM95Zcna+yg8O/Qx2i49GQdc08cU07Kn6U16r0Fl2Z8y0s1robQfrXJ26UX0
UI6eAnE5nu5xIpQpU8rDTwmgtLDT/SQGRpTHlqUq6DtBVkLpCVq2Je/XPtUHZdqHtocQo/CPCOds
yzDwmGPOlxmGP2cIdjm5srbP5r/zbM3aWHlI4BKgLmKwg9C/mjF71In8eJzyfLEKsAjDyzv87Fa1
uJo73GnKERF+RdWwWgeuhtWCgKqYrs6LhcVRsdbqc1A2PUc+NZYDYjcbqMvIePC68WGOqnhQ0Hz3
lSxk6J4K7W0v9CEsmncoSb1mqAlw7dnyXNBktoywQqPuxR8FJ20m5vSk2Q0C7NKs0lceQhiUMg8w
jpPgMUSj1UozAX/bL2JZFvdUHtRDslQJCERkSRlu38WBQEYM/2ojacO4DpLuqEpumpqYc4jff07Y
EKC325yhHeig9nxqWvR6L2JhFIiH/AZ/h8gY5kY+pbmtBhqBo1gXhCK/oN57/VJW+CjuNRBo9zgB
zFUg5LaoA+putjspzL+pY/zQhp/ZLbcli9+ob++L/ckyAt4cdTodVEK25mxE+nKfPtB25uZ5LVTE
XrfkFrKEy5fvWzapimQTUmRSL9RNO/jU6WfbUVsQpFmSvDDbLuwwJDokZNV2DQkDIH3/WELacVCc
1cDNCcxRzuCVBF7WBNhREAXaRRcw0DXcJhtbkN4ELtVbK5GK7zk0H2gq1JSzmsOMiJtd1Hy2+133
Wh0QHVuQistIrcs1zzsz9bxRg6i1UVOBnCrfMb3lkEIX4L/el7SnLQm+WGr/sk3os5wb8yuMFBe3
q9RGWWFzJUGUmtPlLWWJzUNd1hP+cfMglk6atasRiBjo2HBpvuquPEFdANPF058YiJLUAfLy8LVN
qUyQWqF+aF21JBBBRZlZaCk8VsK0cx212f2l5tb5IbreH6PevOViuP7mWN731vaZvO4r2XYLtCP1
S/R7ZfdGGm6LpV09VizeQ61YLsoysDVbFhr9ffmoS4nKmVKoKcavwSxL7UHToBpFwWSPcfSu/QRC
azs0r1LcrQzmjxsBKlSHwv+jWd16kjPzRddysDfq2hPIkSPekJddXPdBhS2bkLTGV064rcH3+iGy
tHUKFMb8zEC8CWzKT4LCeL2yjh2S4Xe4qzkQsii3dhvvKXFgJu37Vsa340X6/3ERwk3/IxuO2oSe
BFcdonwbbQ908qiFVESecRTzjaARGV1yI4a9Ww2lM+MAxq8FYCMeYBYbICpePItS77FJLP1Aj921
pH82tb0vdDOmnmJeH9ZQdxopHDNzN/YjEUtzdAblgrEi2d+KRAJ0gWn0s8J4WAjWt+wPJr7o5Ww8
/SnWVUJaZZwC2Lxo8nrfLNzXGahJxwSV8LBJr3GG2bfOF5w9N01QwU7f67lYvku1o9DtGGlvbDqe
IeSnyQ+cafxOtfK+QT3Fq79f34PARbABQoK7zNjYkq8+5rMpe2IT5TVse6dtpfQRWHrPPziaH2jL
FSnp9Uo6fxDXX9yj3PVJnwgGLlBPjRm/dSkEGA4lIBYRiEjq1qyBEh39x6z9s3Xr1zXk2mhQzuDP
oeXN8C6Enia2v4XY/iOwHF24JylJuzRuM5ieF4jGDIYgVi49syV3weDrzrDJMb0CkHgNa5JjWK0S
BXD2nFZyHc7wjeLTHVjgZcjbKx0SEFVaIWKnB0WCZKnUAOWPzM0no+kksukcp+kM4jvKCbfhsxSd
4KM2+tc6K30YulNpoVOHSTWWaaszuSItxefpV6Ntuh2MbCTJsQ7DmJvUWh/kYv8HDFcDRIdC+Nah
1Cd74uII8e0NvIMwAwU+APpElJejQQQRXuyAZLwd9wHkY4lXVn8qIK61G0x1Ensf7XQGkRivVQ+S
ebhdRXPA8eozotVuRPT3GKIwYkcn7SciYP5E+4uqN0fxyk+lk3wIDP09Mym+xQ8niB7b90AvgymX
6YKbl1IKA1waCCeuHLk477ku1S2sqYfU9BjFjAaJYra1RTyrT6ucRJ1u8WEz2zmnCJZu2xkIYFiR
Kt/+EIh9WFGCmIqdckovjzb2SaUI/POJJGN2SOYAa71DeRfwgx4SwJMTfq8/WRpg2TRi0/6E1zSn
N0aqX7+7r1i7BKRgXX//T0o0JO7NTdKOVKLwj9bikRrSMVuLzrrp6c3oyPWLWqOqsuk5+zciW35i
TGaIvP44w8Or6FZ9kqutF3pnWKDhbTykFe2QlWU4/FsGv5XG0bO1Jzp+EI+4Yn8a/1qtQeFppxPt
9GOD94q9OLU6kZ6/qXcZrX1pS8NBKXmvrO3QhzmVs5YYVgbKkFMZj0D7lpMaxslRplL66WnY95Ga
YhMb4UXToVHX/86K79k6pczNkVOE9V7Dal2mfmqBWjO70POTa1urPqVKDJ3wXo6y5FP5RX9a2GMF
FD7rWMZ7h0E1FKECkEtU9gGvXvbbHpaFg4/WDV1hp65a6rzyCqTg2Y+2K+apxTJLBF/AnTct+Ur4
yt3s+tWdK/2Pshecn4CF5sNfsKggQloAw2YEJ6rk6UYNfCyB7FEcml+5EXhuNpjQryF+qQabxoyK
XE6rB0nUIaYDGhvDuwSGCIBMDaRJP26PBsYW6/D9xqnvVonBCcxJuhAVV/JxDk3mMth1A7lPLWzS
77bCGLmYxgpatS9p0EqFD8FfOs4lMTYFWslLBlwvH3K70jCONOE3EJchRa4voK2XXm2f1w1etEYF
2bOWxOarkGOISCguVVpqWYoPU0l7V+EE70w7BZxnVds71mXmRVHHWxwD8n1YwUNJ+KK0T6avCiiD
mRRttnyRl4TPnYA+yJJkWcmfoJyo0/NyW9xVbihSQT1mVVeh+co84aeFzVt3+vPO197SiqlERsUI
ehbXENh/ue2FKjQWciy4goOtgmcDW0wqCC+qRc1OE0lOKLm6D3E7s/kxAsW4NDi21JYAOGj+so6G
ttXejr7zz/FcM3VDjZEpcxYn6a8EoZZXjCuJHt1pJ5Boc6N0t2MpdEgsGdI6C3NK7MI0QuKKf42+
PxjZ0Lrjm1eZq9R9G1Yo+cvyk4KOSnx2Y7BWCDoHvTLbrvgpZMlsFnH8EZjW+MwOSX0q0LA6PmnJ
Kz4+cPQB593iyeuZzqU1/PT7vUoaaU6P06lYh3TywMglpm+50vT1eAsTLeeKbutUfSkH0AJX/hE3
89MvaaVDrBTNOy3E1e/65tdoGuqxgSc7y153TpUvnsZoQZF3yDTFXi+MT7n1vC6qjxUydVEpWoR7
6c9S2w6Idu6aOoljqOwOzpNJLFyiKw2+xHj8qYo6zuxXIWvkowr/BO7ULf5LWuv/LuHE5WAdxhDO
yNZu/rNJsGPEALjMePXZGpN5cx7RGqe/yWCIeGiZwsewArUE9i16iNP0ahC75WtXZF+KgK2aIh3O
VYallez91mbNDxcoTzcuYWPee8ojmYke6Z2dSeDX+ZPegGVuS9c3p2ZTXNzW5Hj3Sn4Hh96wD7LU
SXieU21h3a78jqnX0FiV6iSfnkjcsKTE1bliM2eYyCe7KgkuD1YjjKPOP/2N5o07aSGww8WjIDB2
IZamHkWATt62l3UhCwcrHORB6sG6GsDFgulsXpPmneOHNI7hx3J5VLLWkpDobp4Sib3CWZrdo5zS
yVuZb4NVDM723KqJiFR2/ld021q6bO10zhfjdB/vnHu4tGJ+IH/5Tf253YJB7h/jinKNya9EkIux
4qwwP2I0HNvZhuxLtcic6yhehs+aM7GgnC9L208eGzHK9SGqlEbZ9q7UKFJMgPGUa6weK7Whe9+e
3qEflNevZ//l1G/HtDbjcFLHw8onxJihdLKlEg45ub1wTh5tQEX2qEj9KSlDY15BDhtWGhnTFfwm
dwN+YuBKgVETgJQoSGWvaeba+JgGx88fm86LawsYIQSuaMZEgwo9pUn22DDoHSTAs4pmzc2qhdN0
AJjgbcI0YwalJSM0FSzqwmPO281Iib2s885dQVuMjJByBzhMPzNMmbfLn+2MowLWT8cxaPkY0zf7
gGyO/0WonQkeLPWFK4tL+H7o3KhoziyjgJtfphF1K0emViDDmDOW9RDqy7xNwQZjBNdW2jIEqJhE
zf0jTflOjrANNPILxBkTLCWvjObEteyzSFvnD8+gECwVegMsjmB8xKeJgbimAcNovQd4J0EQ5HuJ
1KKsmaTtaSNbtjI/3s+qeKFMedF57/q5HMkVmPkp+pasWWugqaqdZjScn33gBmVvirvSUl0lQ/Ok
RVzoHQb6Vq/xxRCuKhmXA+0DFWmLSwvI6avvlW4EGz/3a3ONiWHmDVfvgTkco3uns4riccz/Apjq
N7U6aUV62mzhvTkO8phboB4yYfhZu5koTsia6ehWjKyVYceOR+gKDtNTwtG3bOFlkoTZR8tZjtP7
iOmKOxS63NPaEnYKZrzfLS6LPgeWBZBZ3/icGhoAUXV7Gt+rrnprA30aSbXbgsAmqcwnER1dcP2D
an1rwD7+enFoPOitEUkFQP27/gMZkKaQgYZ1ZQo+kLqr8lHrKPwojbCjumGXh+VZfIlwACmlJaRf
Yl7aXo81F/5Tu7hOqvmKU3RFefSS1jtLPaIxvy3Jix3PDfkGsMxmlS9A3fnsc7Q9iVyOGfmkDEcj
0h+wkQaEIm/3r7vDzob2n48BvFYppdea6lVK2m7TPB8kK1ZUCW8kiJLRU3W23ViSJPBFfp3bybnD
/qKqk42+GGWv2+WzsUXLuXys6lnhoYu0hcPXCI4K7OBj/PbQXoNdOBDOO34hgKNev/FDOlYkcXxL
bpo8unOKsixzi1nJlS9+3sW60kIIWxH1TnZV1LUt0Srf2NQSOocRlrDRDnY3Bj0SUICmO675GH8S
v2DJsOZK5M8uMMyK0d2NUriFOtmTBLURM/MfCcsSNMva6Nm+pDSf8q20akg1uny4xHcaI4/DgTBe
7Y194CXDbkVGTQsBnwFGPks/ORVfeF0lvbzzf9PLt2lgWp1nefSrtafD1v5p4Jeresm5LvB/xNCS
WeOlyuocob5dOMrUZ5tjb3zHoxzhvFuWH/27HKXl+YziLOIcS8Qpy4MWa87St9moHJEFeP0A0BlZ
r3zi0nZbnW4dG1S9QDj/p96YLxZhkUmJRixgfiiDyebhk8DtVES7YPgZW90GdmmPWa6/L8yjdZ5K
9a/f6Jh6GyM0yDLO3RHLW+1I4dor3FBC98BMKw7Y6rakxnjBaGbrbb3hYKrTSEScZxr8sWiAi21K
OKoH6dDT4FzXD07rFWxi7/FW2AAEggp0MP4Q96G9Dl1ccBKEebY2yCmPb0XKnUKtzOI5uu1rxj88
UWDv1n7ymeh1DP+iP3Q3xC/tF6OLcRku+DXcNjKixdvzXN5OSHhXumLJgpOeurgiJBefy7vKbyEA
DRbT/1cDkKgmYRVlpDSy0ZPWOJxo54SgYR9Ju7rIy/J8TtOq7Wp1grUYk4NMABL6vgK+nFaQAqrt
fibLbEXE45WfwXv/m+GsTMATCUuhYx4aGr3ASLx1HVfvUnLZzbIpplKqf04xWXQyeEipYRuWnXsB
f1Q5fMEAocm4q82lANtjP9Z4peu0NWjwbPK94agM6+Q5A/x/Ya+dFm9Fy6QofGPrdYewVXXi+8Gp
mT+UTvOeOoOlolOmmem6K6C9SwpYhNiIkjGFbJiEN8qvUfEaUKp95DNISAUPn7161Jonu8I9N7Sr
npEFZ0J1AaJ3PLi8OIhGtl1yWLlbohAXdRx4Uev1dbdcLjJlmy0Ud4UlLzj3yvS61d1uP1hmggJY
ndLRWABZiym8SC0UQgvPrdg/GEbtCdbHJVO7fiJ8EySg1H+To+eoq7/2Sb4JwBh+3nsKTM2x3FRF
7N8zdyUtwEotRsslVZWvFqlCbRx9TgRBgEevL0uaTaO0c+3LcBCE0Rf2mtIxKRJL8Q9Fg9ynnUGd
PAljqoixIGonmfIfWTao0daSB2w1YaMHYcvCreO2sewPBN6uEkOGxznn4NVe5R+kKXu5D2fgTIS1
LMtrwaiG7G/Xa4V+P72RzGA5k3QHVKM9CAwvZ8vwHGCa5Lf4KoBJ/XHHw4IgZMPQEj2RtYXwAxK0
FpDM7TjoZWIvQQrlb6PEq7rAtXKHuhtqCMC1Pd1ZKVSv303GpDtIHwSiRLaAe9CFzGf3nMHLFZmR
qdvyLzbMO8LA6i15RnB9ZBC0kDSnheNymsbBXvjiQ1CEGcwzGYOE3mgOcnEuMUhXRyPpWo5nprRq
S9Tdg5fCf+xthMx75pol8L+QmiickE+51bfX2kgEBNt5ARZ5ZR02vqxXx629EtK915AwScP2X/cs
DaxzrUZ2ufw00Tavr23BldbzhbOChPol5O4jVBsAsbGS2tWgkXRjHf0R8Y4lybwaB++ln97VDjxY
TkMAfzyBYhqbYXZG1aBBR6jgwphnKHpbVTbGb8AmTiFrLQBmdYfrrtUL29x6onidtzcCbZkj7rjE
zRkOB5z/5DPjQ4IuDgFb8/XIYZMkNqeJxnbke6cJ1KvUYlWY1zqEBH9ITfGBV/xWBQHiMrjsAWwi
sLWOGjSUJxRAC9M9zk2PDygjSWOc7mUo7yVuT/zyW/arTbwdIUsaQWVFvCDYtAHPdj4A9M8YkwYN
GxKNcMjA18vxi5aRz4MXxV7A+T/YKDR1AnTScWzfRBsrP8KzhK7Hz+xlT3w6Vt/8hc5xqteaAD5D
YfS3MpEX1yofcA7Ti2ZAVy1hEURmOZ2ZJsA/40ahVhr8bo2m9Wkxr0UrLDF3yFLlJsy1wR65FEYB
S/BxfBs8NyPJmdKiOwd+nC6uONWdUDpChKnuySLlI9uT4gtpwiB/cNjFh7vxDPUaV5C19Bhp1WRN
ndjr9YhcwmGeOKyZsrflqKgoj6Jfp0XIenZUpXJy0xjURtapa2cB8vePRh+3nZ7uwHclwBj9xflv
ItpYqNzYOoGi1yZRzHZuGFe42eRNJzrbSDtGzbtJaHB/gRjYw1dByBMjIqu1OzyNU5o1BrOV3mlS
F0us2lfLu+XTkDJlmTCVPpKJs2qA09/+pVz9EXnlWRoXdQOvWciz9oUO7e7dEnM83BLjLRjCkmzN
NHKP4TC3XwzdmX9qWSAenwo2w0A+0ioQiSYGpCwp2vrpu5MRbq7Jq7eXby/XcA0Bh1otQZjcGR8P
eMUmB1Xn5DVDO19eFbhkz1pKFfZ/m5MblH8+Pzh2UH1XBjRbPOuJqLs4Px04GtdnVtimh3a1AnGc
1+MoO4tvLbSGI2NwfPmZDzXpZCBcwCeUOY6KAaqJxEuG3Tk2XPHxOqTvvgKg2PJZAPzQfe4FBGjw
i6pxZmDQbFfHXs90uUlt3zaNnAW1CwSSG3uKxEG/iB2SCSA9SUBkHi7xSNkipJ6R9ooBoqIcvINB
H7jMBo4HT3iPXxDnXpalxjxHHaVAyLQ+JSqJ8QrqBE0VGIg1tTUuWn5TD8Lo28psp8vO/2kfRqm/
ZZh4TSrmg1t5Hjme0cKAtWq2vEK6YtSN4vFRhXIygz+YEnG9322jrBJAd/sK84kI+cwB2crI5r8E
EsLEeMW/bACdY6VBP8g1vYNu1lTWEuAYW+Z8D1n/QwOwAlOF42Mqwk6rrnhe0RQcod6PET6ovhMJ
nVZYM0Ao2kR1NtRO5Yl303DM9eQ3ix3CVtirUh3k+mVX+Saiq8iZfVEtGkdMkcOIhIPOZhdSUE5e
eb8nve+FVWc/n0oKTVMGI7Gcunu+qcG4iuxTVoaa82E1W5XPxKWq4Sue6Rg4rmGknQkoGBW79i/e
nFJBTiwnccvpFGpx0oYnZ2Urbrk7XuXbuQVANQ589a8D+a5yex7CYLuwwsRUJuTy73YU9LSSNEoC
XmcAcRAsGZGW66NViZlaVX6jcYx+CFjMQeKpcz7XtyR6fWEz4NBenXjDtXXs3kQm8+1BcqqwQ8Dt
WVdi0VRt/Od6lUKTdMeawpQiw6ozKkWNITEB8gNiTXaSO7Ig1QvGvPupzXOU19PB7/l4EwCuo/db
LExbfmmcluAVGyTRm0++lBQxN+Wyb489ZKANex4+Pa0eR1KcyZgz7FxMCVkKokbFyIw70ghTvmK0
CfB1IXLW2OyMwj0BdDq4kjMMARBfEUF/Gu9DHiAQzdg79MXIkNy6YZ2ZwwMC96u3k2VrgA75Xn+Z
ZBGn1uZ4FVYApKLUPVDo9GKCZdMLqZv4CIRn+ycTLhwjvvCMBtQ9xfFpS6hThKq6RVP4KQz15aY/
YasEOv99qgS4lEnYoSpFa2UKmbbTWbHc5jnBQLULDbVeVVDIxhdTnWcR+77ZpX+bBWQKcWP/6qcP
jMr62tCo5yrDURNN4Hwdw4G1+d2KHQld7cQ3egy2o0G/ZWoAkDTZYeMGwbce9tEjjkhL0sNezCrB
SWwhpAs6BTSX7ZRpxBdatvIq9RbgU7a0L/bYqzcljwZZieLA2hwZM/IcaZUcjbXwE2PibTzKYSp4
gUQQ/vBteOe8ppaYD51/7E8dCi1m/PCprBLuIaMa6hQdtrouOeXXaqMv/I3hi8wOdWxFimiZsUKu
JY8Ld4hxoo9zW/KqkM37G0XIUcgqtibwXLKoITaz+v+58FmJAHXc1UiSPQJY2C72Niwsiw7Hgl+c
WlzQ6688WfDNATdNuEpo17XKdsm27kn/HCWYaB82vr/rEpF9HQ06W6a8+E/ySJcGpKL8/c+sjDGp
Qj2kEpu+CwaXWiKlZ+nAiG57NNqaGcjp/sGeDDuk3Mn45B5AstiO5fsEohkw6VaLem1K5RT1uGtk
WeqoWSxT5P/ZeJi2wMf/kgdmYiNglMLBy7Hoi95k5FEIRHYp1k053L/IW3D1kug5mxP1NfwlSHZ/
j2+Fgh9aZZTF1HBog1RPWhvPK2gC2gv+bB7cwFr97RizIvyG4mbZCn0mqg91wnHGPvCCK30F60mp
nA0qqqebJu1CO+y0ficEZqcU7gujg/G5i5rXq0gsuXg5uF+MazwGtZytEcfPyWy/r2FUk2dV8iC2
TZTMWpK+qrfaBGrGiAAidVushWQG2RdV3myu0PLJid8Xm/cMPXgfIguatz429xuSnTT8lyOXMWn6
fEgNNX4cw0Xn98BVwLrYdErVcfEx1ZYxPCsWhKRaJgWSsWtAisreWwfgFgZ4S5F+FJ0IRgIK0lXn
fs9iovZ3J2n+9wFb2PBbcSE4vvY9c5s+iQgY/rXZvOMdlBtjqcWyZV+iYs+uilN6Qrutw1NZj3IL
KBOaWJM3FUXbhXLtApC2EQh0tpxyKLKfwr08ssu3GM/6HGU/gX4vF6CiZOy2X0u7AB35i0Xb1MRW
ezvAK7WolXJNTQ93OerggPOSSsUKJSPUmG4BFX3XfO5+5fX2Qxrep+KAGnpPTfjaEA0qUYtA2Qjo
OZzcLW1Hej0Az5mux3j2PldCvcYJoLvhTwcsclfA/YJ428qwhEXmPCkzLN2ZYUknHT6Mfe1QUYI4
3jS5EOiBavI9sRYn/orjHbAi7zATX16M8/WOLjkPCgEdE3IbQfsXUowQ3zEkYPhNbzhdeCvSgdS1
92TBwZFEHNmu+Z1lBz5AIxrX/ZqJhxjSx6HoA7v+/nQXcqH9RXs+K10q9FBkKQEyBUWgQK+3LErS
NqjNfmrzz7A61nEGokyiVzWzrfAnNTQ+NOtD1L2OM3JTqfUlYKLsZOG4JS5OizO2dpkbZ4DkSpnE
/an87E/M0dHbK5l44OYqC373wrEDl30Ev3aKP6mz3E9eVIf1MkZAsMwHG9m5NIOVnL11qdXocMCi
epoEKZKuWKaF4IY4FdfMdSik9McuCk74DdbI/g4UyVL7uNBDdO4rZlJimVgvWMnb9LV+Nx4ezp03
QQw7TEQ0A7VVMSOO6xKr6yPC+Gj/S7sOkXh7ohWqndsi9H4v6tBy2BF/HAaCrb3kYi1/jQ1EUuFw
LD9D+42rhOlBqP6rlfvr8oFLzPq5gbHcNTwQx04LEuc9ky+fm2qq60powvY6/XAYl6L5OcE3ylts
SBtFWum+RrfJmYPS/TSmZUYqHi1n/d+1JFHiNhjQZ4+HU6ZpUVwOOfODpS84ZWwYGFg6ETZqd9hQ
08Et/gW1E2leRLLL3tGEnxZF0wCeEy9VrEovQg3f14haWszrrD/voiTeXeKAJ3IdCpoKZYEYLMWX
7mzyNatfpFDSDXOSiTYMv/06JesDWPzn7RnsYA98Tt7VbldLahg94o0enM9OAHpBQiNjG5sJv8Or
DCdj5cWaLhBuQSnQkJYKjz7UBXCgJXbc/bYCukadkxwx6tEqJBaCLdFwJbn1U+4GrkK0RDxwekr6
Sgi7T8BdAQswMks9zzdfqw84TvkRSyonlazPSQU7418ou3TFFoL5hBTRousuX1hCCqXHjdu+mUwY
duiXpk5qPFLEtjCjom4H/P+0icMgYaybqzc2M+eonHlP5zOewsEAJaQ0sp92Hx5u5d4WkTUWsr15
/h5rmZN2thivBgpsySKDwA5El14injjXWjKVLIkNd17B3i4bqzYq3SUkW0Qs67A3p6bZmxAZFrDo
WoFOk3WyGNk89L/xa7Hk03VToFAPEMd9qOnzCSPFhejf9z0gwwKwKsZG2PCsX9Gv3WFbVvPHMlyE
0Z1sL5L2TUnjnBm8/dbvpbMRXp3gkQCDjlbfUyR9uvy9uI5p80NhFkhfnG+ZnwrOvfaBIY+XkTOV
mts+grMv3590cUWPVGaHYRQM16PYjY/n2HFesqCir7Kafer1s+Ko9Pu2DPuAtUaeKDl75guNLcYf
Ro012dd3BTc/hA02o/hiMl1cZ/LBbGPOxDxBrDpZTzJuUK/YvUStpaREYLr3yZFtwxrkvNJmPvv8
PYtvrtmLn4OB/Zy3LuGdDLwvsC7ZoarM3+8yWcBE1NPSHhqXOmtrjvoab/W+UbdBUNQ6i0BDBk+L
r6f3Lei/Bcah0dG9TCW6ZBPesDC3Rn8uDPmgTEI/iDkBe+wovGgrrq2u8u4a0gpmAXV/K2dDzbG0
UYotAp+LliMLfvkNdrpBc9dHp1vtZ4cZqNkUxLQAocIU7i1EhXA0S1MhfhcnI2Ga4u9DOCnVHYMH
VEcqHCtZk2+s1pUIhIk6PZviD8WVnGWHzJW67/vfccBJDC599aWFx1OboXci3qy4X9CeSvcd67Uw
LgjkYiXvpSBpeLhCUwXr97ovyQKgyaKpub2fiRxIG/dHKZP17/9w/qhZIzJ33SHbuq88I/5/gFI4
KHTehh5H66wCK2nocB8y/hRCJxKXc+Ec9u1vvpzwKvpFdUCPfBPEdUmZsM3O6F6kwl/LAe9gBMQx
+Jh3UZns0pN8qPaGVRKGAEmchE9s2EgKAWUCVwg3RhMdV03uW7g86x9q47qniCwvd0spGxLCEiQ7
6Su/BL4StpUqVzsVn5S6qoJPYOvTRdVoB0okIjfHEe2I1nftvE5UeFVr5ZnR7/ZS2BAD6G7ur02u
bWBB11T18sDpAdnsl2Vvg6j2Imh0j5shCX2PvMmJHPrVPsyrzLyx5UUbkJH2LTBgev79Elvb0QB5
g5L05twh7g42pL+nAK9w4sF/GjjLiEGvuDpYfL94E3+0T4ssdukegIukqY++hux+QEtKNEaLnrP0
lzCXWk0O3OPxJkfz7UtKHKds0GnEO5v2JRpMMFD2Ce1qVGlpyJaQhraGXAJf1zKOoY8q4gZ5q3Ju
dY6xeTID2Z0hbSKYD7mrmQavcZ+cJO1qK8XOBMwMwfx+lDSQEo2UGhRmWojkQ/ZhuS2RMJu0li+a
cbg3CUm4nyWRg42UYWp/2rtsc2WO4BkjFwO/n3B3H9ZyVBN1zqV1uoKhLI+LjLlzFRHwHCnKrWMd
/dzOSUBlqXojuOIv7zhBXGR1cZE7/YjUT6VGo+UZ3tpou2Nqp1e9iiUkBPS2J/Ge0C8UcSaiRRDF
NMG7RaQ5GBlSb73vRegEXARAYItMAF++YJJSsBvtcavi3k2V5MIhIh8iXEf+hjpSKpr4RGUAr2x3
UcDnfsMkKT2K71S1CuWxQYfrEFGiS4SE9lPNTDIZzwXmxlTcceYMFaOnDfe03W7VG22Fu80VEOVf
wgufUc/Po0fWs763YvptUPfdaOGuB6KjeP8zK/vRbC58uQlv2Hezaf9UOFITgB5pEBBBTWBP33Xq
eEhUSzU1Urf+How8CIqoZYiqAeQNgOnaMrJkFzr975swo+XgbeYLrXkdS4WhlDn0Cv4s9OdChh4Q
mQuybGkgJyXvguKqa+fd4ZLvHlGLqgh639LpuHiex9D2up34mLSYTarMiA0LU1RQBDjWMvGFsGWl
MV4LhLk5f08odpbskd2qCsDRsPO2Wqtt0JB3M/ILl89U6e1nchs2/1wtLMB4XbgaDQVv1EDAINUG
xLSyoUk9OqeINjb57feHNdsPvPeuaWnRK6oomUoNlWYOOo4Ab2gPxlAriabEybWwVoJCEw5B+x12
V922aorDBmU6vEy6FdZcgAlWtk8SwAQTIdkwXVpP5VbBqpNhgvCtg8gmb22RWKuiE2FScrv1aE2s
LZ45cyRQHE9nE5DWaOWmJ4EqGhnIZmdi1eWX4aEIoHNx0Qjf7AtrJ+P3mkuXcToptg/MWx+hywVC
a92jtvYKwdAoIKbO/4bT/ROWrrdqjvhZSIoBw1hVXyC1vyIHZzB6GFSgZoU77xwyszPn4FjpfBR+
qUvunIM3Fyb2fOiHEVcPe8Vxd5QmvpSIszfqHaDmxwIqoljXm7gylQyo1J+5m2/k/EKyYKuCnlKY
S2663QMipLguoZVKxW0X6PTWXhxi374K3sG/owIs5wQ5QZaHtqJLkSbftmN1tN1N5rCvG9duUg6p
wDIM/eXxO32NEqlgDH81nbKqo8iS7b7KkH6iI7xfDOTimfVjBYeyjAkTV5KAXSM30SMQXnPg5LQr
cMe+G3gj/Ks10Sgi74L8r/0nd4DLyYlNRdzNmgkHb90pUZl/Q3pbqZWe4mTFFEr0q0qx47RPAb/7
HBZ5T0FWBDOm88IraCME5e0RRaYE7b5p7dO9MMJM9aVE8o968Op1q/J+CVj0NoxcMGH2WqAcmM0t
KXfQLQd4vNzjWebxBXKdoaY60ztowOzDPyEr+R1B0NgSyilh9JEKx3ZODfu7B9U+/R46ajEAZL22
QckHNx9hWFbYqhZwvb/bFzoP+cPfdZLnz/8h7ATINfCjGu1o2rcRlpSEuEViLJ6lZavib+dCjCff
BfRbk/K6GOoUD71BYj30tPoAJT4YMYGLiyJ5Y2J7LR2Gif/iUMoLBkVe0mlbDsxD8GAaJN92XAFu
/Lgj85L6MvTjSaaMKMsToNERJXoHyw9NG22B+VE4mszcGr5Mhi9Q3iVTmdXoNOR3eXImH8QAneZ5
TZJS/DeP31R3KX+ypC1R7N4uT+3nCPyqLQMWnLc7IeiPfo96eNEC4mRt1JdBfTShvvFdGnwamnWx
jLWxuK2T4tRZUjOKHKZCFF7CpkFtcUAMGo/YCk1pDqujgj0l0+HyUGWaQ2ziRfxExfMI6vGefFtH
6NlUdkMB6943O22ujN2jvzZHZIpdceYhTcY2ZgD4f5gJWg6qw7OqZRJIJ0efXWyriWkWuNkj+ZBu
sEDXYu0ZOGeQ9XslH68lLjqXXH9zUOy7DylVCEzHo2v6/sEyPyX9GA6P4Lpww3vJWZm1ivBPYg54
LiMUssjSPFMvIhHGyXR1iceTbdUSAHKfWq+S+pRhofjS67MoAmPYXto6ggfno+CDse/Bjg549uAm
0PtdBF93gZDAkVLuzUgTN/2xtAsmJZxLNwBFnAvo3Js73WgJZLf769omciy8m9muQBpNBNxOEZCX
qFkCilIIiL3iYMwbJvjyFWKZSA+wxHtra5tlb2SjYiE5fo3wMQoidDZMFB7bHgHfANC/eP5A/64q
JEMrRKzzUR52xECacQTGA1vmn7q4xzrnahJiVxXAYVWCMt1Ds9Jw5YlWFjHyFbPyNdF+pnKoDbQM
tmxYSCC4PZfl+Egq9ZQ4KZDAXYUn4+yd66i5f6cg/MxWwjoscxJ9SFxhSuMPy3u3+m730C3BQDDi
40rUzrpo6R7eI5oP0S/0hMFngs+A4xW+zLj2OaIJjoSXC2fQZj5aqfzvjLnwFrckKbIImZfDe73J
4hi1WubdaSGYtUd4m15FLO5n+xXrfzkwWEcCYD6v/3tYtFgvQ83bTk00fywwIwqkJpN138LUxrqP
SS/4mtBdbNCnwZ/a9HfgVYgOghcD9yP0zax9KBNAfo8tZJDM0Ff6UEI9CEMXzZpY7C9qSQXODomJ
3FPYAwEm4VVSOUFqfZrfDriXr0CVgtrtFUwZY7meabxY/NZO9Dv5vak6UL1tdD1wUo5dbE5O4th5
iufefYTD8MMX5g/TvW5C1/wuaK1ymfJO47eLGocn7nqiHBE/9Pm+2YSvOwi/bJwzOWne7irue867
j+JoYp6UeGG21tfTezMhXXk4zky3cGSvz3RzKkE8owPwm7ZYYNeNdxVh1pVBwB5wsVXH2/NrzqcE
yyChNvfty2zBpKx87gRUp2f/yQF9qYcWTz/r0ZssTXgcKIZaQSu2qnM83o4pQVOtzzl0vtGXDy+n
ejeqhtft5U9VOJ1qv7B8qpeC2x/V4+BYMlukla6aRcEasTgUfaZyFT+Xd69lXD/D+Irr95sEMVy4
JqE4Qo0/v/f7fhlKI4/akA1txEksFx+ijyWg4mdlLEEAqCgRFj73wnThiZJoSRGN7E4uDW5SM3KX
P3JoN91/cd9dEBkRVQNil/LdCzKE7fIb3Pak2UT6cLclM20hvhPDFBQ4WrEG9717jaYeq5BZrJx/
e1P2xuBoqhHXesJQ8E05SAeLQDZnMilWigT5qyB56LCHYMJzCsgsDZOSGpzmShhH3tAEbwKjptCb
n9D3lHsL/ZXOPWhIxS1Fz++i0UtEspepaki108hbUMuckYoRbDkLBFdk5blLO3t8jIg4OVePdPho
P3QREbXe+veKmOkNRYUZtnIOlF91s10JT1M/M6Qw0uT4qX33+Q4zcuuw0khMi8ceL8I54vSbzVoQ
Ym6RsL1Q/p39tphdZrcuen5pMr51VuiMp9nNE2bnHKLJRcYNW9OxuW7LBVyUkyKMOpqyPlyYSco6
X+aS0S1v6blRuxHHQy8t5U1CfvEKOoMAjtMWSfP9s68Z4Jmu+XEBGwLzuFzVfXBlgSbww/n2B9Uq
7OVXeIKigyPyN//WLv7aJTO0gQlNF80SiQZ5R/fwHJbDr/5Z5SBCT0qg7uygUZMcKjO3gj+H+NQG
m5+jL/ark/LLKUc7fMm8hznYv1WPK/dlgAjNPq8k542qJaqTL9+DCzsFtv/g9tf9LnfEMxxX4OYc
bkPskLzM4W3H5wAbfoLuhgoFHqc5qophzqlxWhNwgz+uHJNQvcqbZxecW8SnWAGt5PKQtve+eS4/
JIk+76xj95knDqrUYhpFiQn9LoTw7TkdXUN5taUq5yJXJ4GmsqrI1ZJJbjfxbgve8VV7D6RTcdEw
CCxF5JQKOhsO3ts0ktdVimcNjHjhgfAwSF1NxEqvGRQR6rX5tsUntWOO2FvJHppgeLfr2MuIa3WL
pLnrkCmvgncKnFL75hbONf2TxgVoifWRwqx8RnxcP9NQo2Jefv0nOqIsLCTlbrN8iovOosqgwA85
H1zJOVbLJL3EzX9P/6FbOULKkDK5wzCgHC2sQN5LWfr2L4NMtSq9giiFSgixtMYkfHdVC37//uuU
ghu4oDgkx5wTqdB4PtSNRsjo2PGvI3wulU/TRentypyrbuuXE0CGIdhjnW0qWZfaFNPDsozF9OUc
Zxb7cdBzdh5QGyXqmow9Y32tvQZ279zVKtoRwHjAubriExmNh78INQrwbWWnSvh+vSnSJTChVqXe
qUK8k3Kc7ocaNTrvX9GL2jwUxXYzgJPQIWOTg81xiw0/X/kqkHuJgD4SgL/BcJhb54i/8YffzHDX
mulH+QskgCAhN2qCS6BINQnkrtRUATYlTzqLBzfQxkZrXwY9bL2zOo8TWvXTNNBeiESun5Ons8RE
aV2QNAeJUnfjZasIwy0JMJ3l13WeT9KemxBij4gglxYJzQZU0Io7JzZRRK6hZve22H9GJA2poQDa
FojpMhdD599MZdrr+ez0Pyq51zVlcjBcr6xptKU7MZ7FDvbrxXIp0Jw4mWwBT4vKGczCpnPEjMkf
1X/GBz4rf2uSutyi6aUIu75DtIXmKxhkJzxVnRnaLLEgWlOFNmjn0WIbsqA7gNpDaEGWCgUZpqD9
v1eZh9ZgFiFEDyjqHQU9TLcKlz+plVuXuNmxQbNLovPyp9EHAzlZAdtQX93w6b1h2Q9k/yBDpWfq
DriXEm2TG9fG1cCBTfPAQc2h2AZYT3i6EUXmQEqQVMDQG6GwpLbDfqbkD/dlGhXLy3QpJtdAwnC8
erVlUSlVXYOS/T5Fcb44Cr1q7+Exk9kMHW1Bv6xEmoKlW/Ppjpwb05lIkNvm3YSIQG79bOrdpvhu
Cwa/nbczvg69/6xL/nFUs8BDjWbCjlVavOHM0Q30eEfDiloxamyz3wp86zHcFS6xPx6CqqUHvM0q
tcZnxE/H1sSjc8uSBpX/lhIzdsGzH/oOjYNOTkBTqXLnCJ1rCLN3YTvMkZ28TxU3DmDvR/6wYWBX
lRkYa1XDXrsgKAmUHpIjv0REKte0YngDImC+wCWaExqi3A3JmhpNIBSI9CHp+CdXheGGd2r/5633
Pwq0zbujwAIvcVY400vylUHFsq3jwML5ul+N6DzonsAm6QraFYUYRzPy/sRN2yagq74FtwVNVea1
L6suSBi2FGYFuQLE41hXIdDnKjZf5phban2/bC3mbRRZamec3jhc9xd7CCuCYloXBDj4ZDtjP2Li
GkHcsQ47OV9AiyDi/NgEKENzSeAjJtOM8v3aLXfrAfsqSFPbZIfe9WWpQ7qZbO7EUBCTBKWx1rWA
EO/Ij9ELObAH44agT+I18YXErwwepqYaLrVcJEAyVL5w7xz8pYiWjJj4Eva1zVtAvKkkcLsJr/IZ
UOJMNQv/horhnA36UNx3eN5DxH1s192rh8DD2Q72ECQV8/OCwfongJLXZ1EQCd8RrFU6Oz/UKKUm
ntJGAs7q+m0XJDTknwpXdXwPcPZU3C9vB7buuPgpdWwe9lKRHC+ovG8wEzb0aD/AJHGGFAU8uSDI
xjOAqjTeNJ7HylnVOxGGzhMkiCOw72kiTelm/W5mKwgeqFoUvrZTsyyaSjsHur3TJYUWklUVaOXu
Dtnm2f7dta64AhYBbDAhbsHRqjSGLpoFEjy0wsZhcstH8KSaZCTGrxu/SYlZeL28hRUX9C2J1WsL
/kAXj9cbRstiaAJs6oJbKn5Q+JdpxukNaSo9bcF1c4iJJSWl0nZdT0FFSYCH3gt0Cjh4JWblSPId
KLJ5KLrRDbjeXe7xko/e3Nl7KRO4FXVtB5CcPhu0pcFOmFJ6BnuJWYNSc9PQCROdBCac8ACH0fA4
XBIzL5FNkRvOiAEb2eOdV2hBQaEkfMHD9p5vL9367QQdgIrUSw2ylcpMe+tTQhv8skDmvUblrvuo
onhvgLtUpzQbkwXVsOSi7wnnd14wEeeGus4JCGFn4aEcpX4j6UR3sGm78oif3CbAsMLiRSLgoa9F
nb/rWMXAw0VwQ5PVugKmZQ0Dro1rOhEU0Y/+rrqLAhUksOW3fQMZDbbkextcJ/SydQQywKF0sQkB
JjXARgD+lBdcJgfe9E3ItgiyQJgACedlRoWs+XJNWJ5aaTszlsv7IRHp1P5o5eThs0X3BKyVjTgR
f/5X/vEuKr3DAUf3LXpSIJz7dsKoLjdxkwfa6KC4wWA4BmuT+H+addmbfNNP2LXn5cl9m6CVg1JY
bHM2KTSaSeyq9j6W4TqFpebksv9PkghN+YyJQZ+mfjTP751foXgB6p1+6Xcw4pCdE22aSyrhHFx7
sjyjXVwP4cB82bD5TGGPTfj58WWoL4Y5pNT4m9S8fA7m21ZkCPrlKSsOhXp5uVV7yyuqXwTaju4P
SWFGVQMJu+pyEMVp6gyq11P//tHrJ4l0W72P36HU7valwrNNPFk3G0mqinIcF26baE2TrYbwfdU+
A/eAL/LT8DgBBHpdU7+pXdLW7J7JobK0tfJP81gWJOMgVW6QkSNhkB3QXAmTzhbMg1rq5WiXhQ8n
4K2MJiGzPug2OBkJksK874lFWQ4Vjti0XM2g4DnlP3VrQnw7jDrW9q9r0/NhhRWmFeMZtrY/dcdM
95JwYas9XItwraAHroW5sb1xph1WAMbwX3bLIlvhw1QFari4m7IuKIWSuxy7ZfOfuWD9m3wFe3rQ
LKeLhCrOE3spoRZu2tdHWl4WRP0qVujy6VCRT/Z2Sr2XH6VwQO5GruuyQ1xvnclfhGTDW+l+wqjX
lPoLmz0Sx7n1RVKt7ODTFXcBtlwJWMwBAlxXQbzky67f+Y/Bk1htD4Uoi37UCeAWgcJTRCIUbO8O
Y7If+AJm7PDWuoWMNabIHbnL0ljgD/zLWSy5Cb/56zKPwe5nFCGiSw25lGOfX06YscuA7GlDYPXw
VB+eeehevOZsANao5d7jPXKNoIpfEpuBbVFKmapnxWR1XDr27EXtXtxDy/37eOzc4+CwTU4vXeuF
X685Hc6aimaFiuElTZzdB5m3jAt9KXNH5sKhoppbrDywuyaIWNY6YIpRKdAvwkpw0ShOVVpeZzHW
M5KVBx5bvxmsOG3eB4lMHFUwg2w1jtT59a+9xnFPM5p2I7/2uw+syaKB/4+V2iL42hhru4owDdU9
rrjJOtFpLif+tGPfqc0b265HHZDnq0hB5Gn4QgM+PYwW8p4yXt6qA3crcxCDCzQg1+MYAYUVUHlb
7K/MfccJi28Gh5zYyVbREeksYGjElDklbj9jlWTB5CHnzAjhuGPsq79U7Gh5HMxO2uLW1te9F2Bv
6rsvsx77DDqvqIybL/smho6OhxbpbeZ9E2zlSVUjAmfiQxWlaXErEonMwmM/dA/avvuhKN1lRlXa
ClgAVfWPA0sFTLN7z8CQscJojE9oiY2HnBcMoaucdnnYfQBhJHagVEOsFoFisaJHiDMe7SOT1MJI
rm0lyAWmKnhx2Ew7rFIjlq8QY83Z2QseCIA+sQ3MxrsI9yOa1KMRqG+jpkHEi41sP5lApQqIQB0i
L9PLfbLdqg+qFE91ypM1noy01CCEvHOx/YKqb8mVy4VHo2k5F0zXWqKDK0tZ9qDe5T6dn4cVO1W1
4DDrAWIi4wzmFLMzb3wt0gs7x8wcSfhmtDDWNmk3SwZ6NsVYeNyz7KtqF5UeSu51biAMioWN1Lwm
WP5Z1WUoxxAK2VZq0m06Uzb1Mx8f+shhv7QSRH+PrpjIIZrMmP3nGdvNlA/ppFpoPoEQi4IbA3/i
VeZHKv+/ob6lF+tSRanW8F+B0bdjzpdeAtESLZ1aFM/NmgbFc8PsnrTIhnX9VOeqkKUARsdWtrXB
s7c0AG/A4Lk0cCZhAqgA++Ml3AzYGjJH9vDnReSX/ObsJoN6O6a5acybSBX0RSzCIGH7wCUKvypn
Gk2eDyomXiW3sMHZKWE2FbqHdZi4XkvNX+xS5qqqK4W3bqyFCouRUpFbuanlmrwvBe5HaOLUxwWc
xCRdEZEgaeRqqcpsSICEQIRRkHU2qUhkw4CldENEnpKhbTRHESm/i4F3/N9z81m1ni+G7P1Znqtf
TOqa7OzRVaaB+He2LnegjEhoF6HFDyI/GmCwop/EWpp3/A6bbNPA9+YR5EUGvDLzti4Lo9WPO2tW
Ho7sevtGXCBJ4JbIR59C8OKksW3eE6kx2ILcz3R6AkRH9k5VSBJ2r0bfDRvZVrZQ1q6PiuJpLurD
GuvDofZX5awdd//pW+yoBjhZFyZK5KiXyHxBZ4PsjtUlkuZ10v+O99gLHjEPrTkMZmhrv7kIFcpX
trgdzverWEdTAUHfquZptSWYYWFSXnyJDspe7aGKLSqrcTqvCoDUgbFySlhEcXno3DhnfYhZoO1a
T4r2b49Vf6UD8MRHMIrj1lLWRu8fHrdC1T3HDz73T0KwNwtdjB63GkO96cL/tBTOPJJLURkSy+yV
T3vtg4iYsfHqi1/+BcCLvr8OGGesHtRZDt8hXoVf2w3e+9TOmjFErMaKcSTLbX2ZpWJk+kKZjO03
CH58O1VUad1jPXqI8Ulugt7b72uFeHG6CTgpWvQ6nvAOZCJoEHKdc28sgjbFqi/oSD6uyc0Nha2J
LGZJoQZ1bINPcF1Bvqd1X03aHI9DoLyohuOkpmqAW/00oL/Zx+kZ7BJ+oIAYqGMWXgPblTiJFr2k
FWVf2z73HjkhK8ptQ86bYmk9OUGDHaSV4rCRnrKF7hlNWz3I0YeATROzRYeLc5hZhyaGawrdJpgz
CT3AV4uWqg3KailqRuMvO7+n59kkWyx9rv5qsFDWdAiQNJyfUUK4wjcg5xl/UpApTcfomOq6JLBQ
K0VquPimbeMrO3RQie8MJdPZHM5ky3YgzBlE5zO+s0w/2BYVI+BGyIiODbeacFj36hbgH5D+r1aZ
HeAMYYB6cmYEyfDtZMpCP50Gk3xbXmmFVeEb2DI8YRDDO3ueMBRtRrDDZ2UlxGFHnAAMz2h8tKLj
hrLfz8AdOT0eyy8AzfBcm3dMz4cWyBwcVPSeNll9FHeye/uSbxAr6V8fOi+lKDRjPyFAbEXsphuT
HtNzVoXsksJL2+IOszYSj4qPt/6ppB2Hi+up8cauzsZb8fMC4qknMOWiCwzU0QKr+bdfVAdnScBe
NOgcNbef9g0ndkE19fLEnCaAvQGhjEJpBtIUiYMyOt6DkH/ppIaWrPzUHZ0qxpYFifw3/4CZSVuV
ovajH3ZvFMNkMVad95N8wsEkYFt8S1/KmSS4RkZtNq7C3U7jXfLjKPg/xe4dUJXXS71nkfGxqLc8
MWjgAm/D5tkpP9HDhBcDR31UiS0fwvmjWwhfPkqNIG8+S5AEQd9E5hH0k0bWSeEPYPBxAKPb2Csm
7hbGMXIIHEn764Pkh/1aog83IkUagZ+Boju5pI7l8J5ao3DOUhLEouyRWfMXzDaaNn4peWKNorpt
pAK5cLS6BhgrhfFGoStHYEy9EGPfqfRDqIuMU2w9B7o5O0CwDLI+FPomri0q7pKIQQ31/iXq4H/W
NS3/qIA5iEc3PNti71BOBX3qxENKwz0TRkMizYZ0h99AmPGpbP74345sSh29a9d5WQbLHBvXNlix
DW6XZzSuCb8eKDxaBE9BwKPQDH/VbvjVcdis+xq466hfJ8djWX5nqv2hTZM6JDkXI40ZOdIWW04W
34ClGIzJbzrk9nqfuCoaY/Owlr2C2Cwo2O7SHaok2/81Sjk0XkWlaKds4LRYrDZnfhmNTZWYM4ql
JG3TlRxf4Hm966dnK8tLqTUCD1k2hjRizi/lJOZJQYYBwOXOBYwjroeH15PQxZzUJK+dlI9DoPxy
+xtpsUTeVtF41Lv41dicxD0vs/vqF3k3auXUA76EFm+oqQi0MdtyZt1no4kKMFRNbwNIhfWzbz1z
UzPgcB4mxKjBpD8T4fEryklOEnjJ1hDv72ju6aNoI3N/DCAXzW2Wa2ZG5czedE2hwftDnIBhhHzD
75nWSdYWF9AuCpu0HQTfKfQ6G0vzbEmNTbWvZ6FsYvTBc/LZkrW/8ycwVpUPEs24ntfWM4owD7GN
Rww3d50bV4skUXdymHPv50XL3nRhKCdCas5tM/iX+lG+vxlC+zUIBplxeU2fRMjld9E2On8Ikzup
qD2PQsJrpESODhyXeVsRi86uWell3LIAwPnyElCnOs4jC9RwJ3i3AObm8epVHuYpyt106WBO8nNS
plW8ju3WQ4o7a7NtDUHZgSVUDy8Zo648VOOs0jpvjC4aeo270YZp6kKCli7MIKBCdBJZyTJuGSZ8
Ee2v1NfrBaIc87IZEhdFqHGCBV2UZOMK28jPVEU8OkiI27C49drdl1U2JzofzKYlwXB4v189kpiY
+wiNZyVjtFPsmjZQRjoFFVq5wv7G9P9ULSZ4ys283bXwku2e91BUdJzGk9pf6K+LTeBPBOY4QB2Q
xMw/1fzxmWMXsfso+21fBsp3oxrL5E9AVwpKPvSxdvBYHg+G3RX/gXzHo7v9J7xiFqx0VCrhyb+O
VRfMkgQVKsSMe4QSSSkXmYJ+wW0d0OZkc3V6bT17LDqQiMK60lBIrKZjfua4KzOAXH5srvqCpohx
Ojn5/Zx1CI1AW6E6rzhSjnb9C1C6yB2ioyjImUg+8hPT36KEFxW4PHwJP2sIfzx59cC4JAtQJide
x/J6qiV7TPb205GDWOQl7YzkxrqLB+fPdq1rSz3Xnd+U0xQG2ZGjZPDiVMbmxLQfHg0O9Kw4WcHH
H7p6BwXt2M1zAMIW3sgNBpYlzH2HOQGweHBuBKdfu+yn77vaBIIkuJkF6FUwoIXFZ0EAAJr1dann
R5aLWDKdMPy9I/13G3A888wSccxjrUqsPy2+rMp0sVvil2cmF3waXLEN+I/MxNWNJE3k8kSPMtIp
zNkaL0k/iSKBbjVdFllk6o4MWwN0UZT8HIuuJ9qzA37pBjekNz64LnNHBb1OIxx4Kxq2t6B46UBD
m3TVbE3MpEa1qwZ/mCXg8xNO1AdYs58eYYdqQqijUwcJKqdnfgPZCzOoAWFuOmFRZs3cTUjyc6SD
1LXrk35NVBoFu0PMrgOwb9aP7glDFv8gJ4kJACe3WN+gH20m7t+qxkyd9ILA/M6JpF7dItlCnn5O
byih2OL2jnPLY5c/3GOzvcM3mjOrf+WwKlTz2SIz2cJCwnunZbOQXGbRXi8OUWtRlMS7Wvx+cahS
d5X/2nQ6Sd4wHacGdTQg9YRKwfQLE4r1ocXcCGPqPsu5VrB9IunbZH6vch+ENwh1KswfWxvtRJ/K
RSH7ufkTJMEcjUyD2KE9oz2QwMUuprFrP+IRlqgcZDBea7J+5X9xv6FJ2nyxBoh+N+5pl793sp5n
bzArQ6dwK5StLNy2qYA8S9pLSGiwwS3nu8nFyMKQ8q1Yz4GTsPt4NxxxkudIfu8fJdgnhnT+8A5K
KLpYBE6SPyBLYks36J8rfxeO5WtsLQKAL/TpPcz2sHVBvyJOo1R7M9Wv2xCwAiOtthPC85D0XzcH
3NKbqx7YE6W3nU15g083AOqnWW0BkJBKAx1i1OQbRBFLexaqoklI7GWYipcCU7kaUjbTeVeAPilI
4odc+Ze+X7Wq9uLkMZsLeHAV7RZGgbikJ9HpbDKJuHaVLGXDwNgpHwyJAk9HviKVZdtbU/u8QuBe
hmC68qsSJElzwHuLsbjsczuW1oMGc602G8p6fbMqDTZi99JjyCfMfc9EUDOJK+yrBQ2jrGh/DT5z
aG/A8ZV0LgVQZ+1onUKv/CLS555jctRUfxi5FDNftpwCERGxX655/Hcz5zx2Mir2tQLEhhRG5AKi
CVFJGakuvb0Ub3MG3/+UXAfJE0VBAg4yocaEtfl6apoJXDCM71GYFqESifo5/0IFxcYbJAA5xsA0
2rzXh3JAvfa4Pjmbz5rYswH5XPs6oas1xiAI10kUz/MH8rwTDSXyQI3t8tPZoV1m1iEABB1eGthG
xB4XbMimffuYtdM1hM6rPKsgo9BCXnK6DBrpAkvmbZgJYvP/RtqxXXE5EvNjNS8fFgk+SCOZqsZi
D+rOPtOOHrDNWcZTBjS7gj/ZCg79+sSQJMZYmcAjyW7JsQwH7N0Mgc83B1o5GMFLhc6CgH26MO40
K0KOfyP361OONYfAz4LOF3GLxR6ChBa/iBk84LtzZCx8x0syJ2FybSh0w+W066ywmOtRK4jROgyK
WJZ/Mf8GpeZzip25nN3QinHRFv2OUum2+DYP35LtYeHGV51Y9wJzFeI80L7mM4nwimEZWZKRoLZv
/3gcvrfvKtDVZ9i0/DFPQrMFIyVuQUv/GtGhAZTBpm6CWk1Kbp8KPwwqMyJlWPPAFGmf8yKStwS5
oGoHn1rL/u+NlYJjeSxnxBTKSMZur6rSqpLDZtG9UUT5gxhZDVh4QUq/HZ70+pNBL9Fot0cV+FcG
JJba/2oubXYsspzKMlwa+feQoFccs5mRCU42hyP9kjkew3uOVVULrQr/LG6btcBlRSQvuJHXkDRr
CVTeR89NTWHezdXcB61I7XWggWmkYh6VTyS6ZTdHSQT0zlo2ZDRjFKrKmEe4SqXTITpfBdVlE8yJ
z7VV+GRQCMSeYmTzb/DQnGEJp8wy1c/yk/DRyhNLierGac9cL91bmrnemuR0AAlZJ8WQgQWEe2++
c0+ypGjq/oB/pzuBJ5TlY1QO8xHjvE02TmdIzaMnVnk2DAn+7pBr2VF3q2FrocAWYFNy32RSaSiM
2/QitAwkUd0GBQ5tNaMRignfOrxjGMbETgHumZCM87LtWpnBMcsrtu0cq0207aTpBSz/7aKltCYA
PeNDcykPOMGLwZbm3gdt3SVX5WRC68IopQWnZAboZJxiCm4RtJjpCjKUU/QGCuNyXcQkxkbf1oHf
eANtTaviQyVOkxn57orX5J93WiAfUBu+ejbmQHL2wsW47SdKuaehHfjyoSuTuDi7L4bmfT4hBvgw
LXCkLGOzrHBTfam4++k4MAN31/Mg7JpyCnRouCiALl+Xwoxs2nnTfWKHFkltL7vcZ/UydaHQcCWu
FRt6gU6tcDsu4ElwFZ1ID6PbGEzir15SL15BJdgtDJAuEQBMBQGY8/rHSQG25EzMWyRJ5cqZfBWf
P7PH6SxLNdvwRi2v88KPA0PO9Yeu7JZdCkj1Bwr2/AjVroN9Poceh8mVeVRwFphRccZEflmUg0lu
Q6bG6xsls/5ospSbFrKlZVjnZWbCl+gJKniLL/UutHue6JARuxGGAiH7vWDt8fL61V4POy6ojPls
Rzfxc0Wh63Ce+4VWsqcfgzWWo20YFANiHvA2tDaeN2m4hHh0IBTb6Q+62g9J9C9ANNS8PhJQc3Ky
MqIDjU3PtTgnpNIvabyb5IfujvBY88kOND2GVjrxXAU81pT4P+t4g2kFQt9KBC3V5nch80sDzFQQ
oELe/LzokDaaZFAQ9LIYwwXhcqjQsv5bH7npyBkTUIYfKR6DkNFODRqxAjpdIU1NWclFTHJMSGNX
yXrkjRrbppa78lmpCZo14/DLKEncdV3lO2QpmpSmloplw12RTsesDgDBkg+lp23RE9VV8avcdRI7
soFW94Y/WBsI+Nyfl3DrDre+cG0qaiPPUNiMHzbxJV4lzrB/nqPZoel8JPF+O4PbfP5hqR6tsXvJ
B6f0Hi6OnfXeNdwEBC8t4V3J/nPNWBC38Eo9+eFwz1TMYO5ejgOIJ8FuAEXqLBIvRQHm1LWjYXuK
+RcJLTT+sfpe2FWmiZ7bP1pKkgiYAkn2h3IPdslm6pKeGIw+X+5k7/vyz6fv8x19fc9bLKUMwyfE
vkPM2+JqJ9NiRUrUXlqVOzsPtmf75pIyM77pOJ5OLYdAkwr2mO6uVOVksz8aIOVE5zMUNIekmnI5
KvANobsEwpdvyi72LjR/vxvLQijH6GD1fO4HbxIvQw/NrCirPerAhh/pwtT+EJxXO35waRLyZglY
x+n24Zing6vKSDf2tQISUc4r3YoBW7BjYSn9zPNnJYG8gU91qNAYBpIuFHf/Af4L3L8i1OV4eVry
xo4Z9jsLzBuphv14CkWm+5NpaRJjp8VRdqN/xyu/Inx9B3XTBgT4iZJT0JDK4X0SUyVZIRFqOj+0
0LnBLRkTwYi7a71h/WCDfStpmBHSFDxwWJPIAKfNbeMcFpb3Py/swWMlnuvO/KdP4Lh8ngnrvVIr
VbJBYq6IBd/Cs9h0LzR0t5qwBJJWpy8ZMXUHXvd2NWfh9jKGfGdop6umSVJDf6/cC3QIzSO4PWTt
2Azled6tCVsxl1a2VqBboz4H1RsBF/PKISjOTouTHeValr5oQB+PhcmaZioQjT3ZfNR04TUjWJh7
o2QdM4JXGJZmQ+xD+y2kFREpRd0a1mEOP6gZ3fEIZvZ+OVvqHtB9tXZbL+ZVoeDyvccwKKpGSbkP
lHKAgfc1rArsuNiitlxqBEUTOG9a7k1mP1boGAb/qfCQglCpn4016MW2dbrWGA1D0biop5/DDeJd
kdSR7kOdw2UCsN8awXSNyIdYAhVEYK5W6g3TEaHSO0CmeVQjICVNCP2M0OnTEQ8VQzaHBL3GGRz1
ByaGLqSEu4MJmbj1Prkv3+kFgA/GUXgzYVcQkEMzDG/qvID1JbVDGOHb7+KV3w3xeWatWbRa7OCm
dB6rNMH1ze9hnrik6HLD/h4DClvbBktptWzyHVxMFSSdBS0+c6knlZuP5sT+UzFKqHs1sWCTBtJE
TQwDkV75LyV2kKavX3xNQlsdrcGWz7t2yp5OcVAauauU8n9Kj6YI0tzTCtLbZge/NESMsxYii8SQ
lH4F9W2I4n/DsT2PZOmldgLXhEqrLNG0o/rVV3CDiDpjkOeKlGj4eLBXX8QChKB9RvQG3ZNFl8Ti
9uJMTyYyawk+wf/v2D+02ialbS8siodgDkwzEqDAarfA96mVCCY8+VpY+40V8Xw0tQxZaDejlegE
SBFznMSbqfqCq2Z/fmOMGiMjayKTLUK8SSMGcYKntS8DLJDp6xvxKAD6taNhspoyi+sytNfGGR+h
/ULokCL5opa73KiCu+CRMuLwDLktrKO9XVorqtST/AbsECOVHWEPR44u9I36Freo74SSEFNdwr5s
FcGjWiNMHaPlXTYotCMYC0XBgh7XDVxUl1yRtlW1kg4LXfqf0eEOGg8LW5sQT+SqjxlJpcaTvkPq
BqkvOD9VTxVG1tyK557SK+2i+0ihBQuJaMBSnXva3KiFjKOsMj3/A5r+ENGq8lZdXlH1P6vVI0g1
IH7D4iCxqo3OvZGUZcICVEMrX7G5IbTnYGY8caacxwLg3w1LxiMDhhgUWcCGfR5kNvcsV7w9c3iQ
JCwIurhLunIhE6awEmg1CIe5emX1DZbcnfpx6azNBDxhlAwz7J4DA3Zj0YUuIDUPTEut0EW+3lL9
2PwAQ49gwRfvHsTjb0hx14JEwmVEevCzUha2tCXK7G56WUXlyh9TiZFpffiyGcmmGCCeiGxKJvej
0d5Ij/lhwBVraPjICF68KPKgUDML6S7/mFblQFNvZLTm8Sqce5kdzI3SGzyzKaJ454hl2yVdBPoI
h5IFcvEUY/08VIkRKWGFFHz4c31lL7yGIbr2hivL6Rl/ZLvYixWfseoUWiAtOwZZkUJ5JH+uxGfN
TLrQTgcH/Vg7l9vyWlSNTDv8gUzD+xO0NeSJnJ522swwglN8t9LgqvNUo/erUW8uWBDCu7PAerA4
n037LZzBwYevVuMpohj4jjxfr9+oh0QMzux/M72NNooofrYg10qiwzzv5i0IlBAsZVOibCYxddq/
jUbiSXHfo4AO0Npr4rc+ThgOPVqom4RtCa4RGbCuqHZfunEN0Zsnv9/1FGNfV/p0t+r1Yr4uaVCa
/17TMGdgUiTVdZiYEht9jQ2/0MNYtD/Rk01VXPSbI8w0qn2TaWIrVSEq2qD8sqK9eDNFsJyqVrBL
IPzX/PGGDZ5Vgq8/m2E8Al8z4wUcsP1k5ocr6yvGSAHeLUzX/GR5ww+kzPRv964EP08iGlVaNlP5
0/Ug2HUwgZTrgLRokvpwJrgeUMF++DCtyIUh31nPeJhB88hlYpf9yHQEWq0VJQfR+amqy5j+lVqV
XtmuezZhwPqO6aRy4hrp9z8o73Se4UrM+LkcyWIL/Knm68rJHACV4PcbAGa2qSa/FIvCnIHRxXjJ
Kc6FVOFOdhNba+P7tAZtHyCVl3SLbsYhRnfS0vfenYSRShMRWGeg2Wxq8nAr7k7eLaFPmNWXgu6b
aOczdvemsu/959Hjj+HruxVNmq50kHkGthGMpyVpYgsoPe8mndXJTa5Rkrjed4VVbl6AUsPoil9+
qymOJDYDr/2B92tm6bT3Q/iXYsrwzLgzErg/0MEdpUKVxACOH+nSSTX799X6IRq01Ch7zt7xPO5S
9J2OzEmLksZAlypCM5bXrZESO4MTeO8sKjwFUFerJGet2GhOsa2l8q4z/NokUPm44fY5GLJRlg3W
DGBlbZKCFFH/nAUxCpLq+/VESd5Nq51oALkzwY+gf6NfjM2XlUOV9FJ8ZWWX4gETEk6PdUYINmPX
lUT7RZMiIIjQzgw6QbNJEU4vKOF5otkmdSHPJ8OJTMc9010o1HUkDzOLLPRkOxMT90mea5DI2KvY
hk/lJMBGF6QSDjxobjB5/9XjvjuNPsl7WHT93l2ZA78Noebms2G1bWzckrhUcxYuTfRTIAwK4VCp
MoQ3edIW0jxcWqkVFo3nAAVmcZ1QQQ+Al64kv6B2N356afRCA1Lms8zSvSOSx69+1+K8Zyuw+3p9
ktH3jZZhVO3szm3iXw1rutbCrYr+n715N7YeXP6qNRIMhtIC/Zn4+b+qvRNLMeCYJCVYgf64RPLE
WL6XD7sajGUJzIrDUjbpgn1N3ZHy/iGBNfcnn+2Wj2kqE4ggF/lpJFpfWr5G51mUcL/o2mT1YR9c
34zMAmWkX7XhhlA/3PoJugNnXqs7o7r7e8Vgkumop9hFZ2h5yOuKhBbMTY6zt+1tIqVcQwZohBhL
9aKPhgHq2pen+AmI6rigE3+dtlylGmE8WDuabDFnDxPFYveYAdZp/1+XiW6CDIMHU7wrNmPxp6KD
zFfsiH5h2ZD8U+AS881m81P4KmNqgc4sKutG+NHiS56LtB5J4ErrChobkb6CbTH22LUZxeuW2d5G
hW5yDyCf2vsHpIr2yGViCbZrcy/VkHtsROR1C45DPawhTPG/gTejWQ4dsBrn509fy5XJium2FGbU
AkHMi64Q9trG9F+gKkQpxI7TBFHCEsnhGmZhns2cb88Tn3+k+JSII/1iW3BMqFiwhk1gbxZLnPmJ
HavW2ZJmhoECDRrr7UxWupnRI8kqtAuweAQqfQBE7vXq9PmF7+5smBo+aoCezoVQTsvM5lpaoB8h
8yaGvXCU+e3wEVf34YdwEBm/mr22MqMW0s8OuUycEHvTPJJVCjmBr3mPQQOAw4AO7awxsk0LgI+b
0BxxlQJwqEX925zd+jRwN/7FbZ+5BylAKWiniHuDC1XEZbNHkGaJdAu6reeF0NbypnYaChmgquGz
7b9Rw9kQiFk2w5e6OZPcam0TWwjymqvlV6GNn4NUG9nAB3mIxsB1Irh0wkFo86qiYdhbOOTwAZ/N
JepM1BUhgIodEA0CMmtyPeX6qF5UQ+1CYlT05qvkmVOE79O/CKzdPlFpkDKLm/HF01855Eo8Wr6c
yyCr4rMvD8MLdVAwANqNtHVmRl4tQDLfkDWlsj8hl7T48RZREnG+zQwVj+0FePRRQlD7o+iAX2Fc
VVIdsO1DHFcRxu2CQcRianIemZjBS6F1sQCeu63wb38RDJcIH4zHqwW+hPf2x1UNMgpVez6WO0+k
UtHLYLMM3K3SBY85Od8qnMJelneBbrL9Gbb/ghAwBf5MrfkX+VJ8vkYUms5p3qJdNb4z930z3I2i
kolsivKHZFPh4gXs95LTo7iv8tiXdqbKOKU9tmZC4wtDP3WFL12uHJd9LqdoH5E5OR0XT7wmf29n
W/Tlt/7O4yKrhXGnStjj9Cn1xbyLTQKlsOTqnz8q01kW4YyuiVMMIQzBDmK82h6j/f2hKcQIyMAh
uuL5g8nyj32Khb8FfB9AjlApYbr+f6lmWSry/4YY5G/z5w/zUrU8KSIq17ry0tSye5bgG9YctSz8
jSqcz4/PUBEquNs2ecydl6dmotf4t2tmetb0iE2dpCyY5mxB9unWXKv+LBa7GN+/dy1279ukEPsY
DI9aHrsNiYhei8/YPCbFuE08U6Dlndgp/LsLzGlTpC/uoNlnvUi3i1ekA7Z6IIwzwRqR0IqPSRdT
USxUl4IPjXaOY00V/F4fX5DRajXR8xWCPLBs0t8NdG18gwAOQVcH9ZPppfAKm2iaHn29lcqOm2di
kX2yJeixbCiCq2OM+yqNmSo5kOR9zNfEXihxD2OR/9JCRKgmjCq5LFYCM82IQdxSCmFVFooEx3KE
ZN3gdJKrR7YcRbOf2tGy+8w2X+W1xjYDbF7vQREWm5JL38rBd+/pGPokmGzBHoTFeOUtrVgGGF2u
OWIBopa1M1t5e1aHW6AOKHxeuIOYskz01e7MkKFj7ZiIZ40A3hqdx/W8eiSYomzG+gco6I2fHBJW
Xs35ETETAhpQK+cP+3+kcNhkGEyazuy3qwKKVpzNw1NvE/YVXFKwLrs6S7URphQmZrK6qDMFLh6+
wmVtN8lQpTbaYhjYHU9QbftzGbT8S+1eMW/4nC6kpATPXzIVjQo7mHc8f+29hKOJwuDcco4rYczY
q9xJgk5gDIEWLatoY4sMKCVMzunsXQ6fEjoMjcmZsZLGC70HMnrwD9MhOu1kNc47mTjpB4oKBoX9
xK4id3tD8duOQapjfQHHkBAyS4eo1mAAUxdKjm+JDSVd3QFgSIAzRJlDK1lTwT90uE/P+x3l0tca
jTNZCF0gbhijswvFBNM05dIbhAdQsL4SXB/V/p+djNBbEuvBNGzTiuvd57/NOMXbwc/hNh+XuS3h
uO2UgyU/+2z3GuE78PBtli37YrcpCdTBK7qyZrvqKs8TBipPgDJKnwTDQlS/nTyKM9iEBb5a8EZe
AuwOOAh+/Lu7dM0vJcJYRTCDFbDFejTuJXKgQdJOnW0e/l/v1jvlpa5fd4IHUMvixId5rUx5uBft
uLbX7RQ0DD1K1oefquFdNlWDBn8NNt8PjeS8Cq/I2/xLm5LYN96ZxcWBZyic6fDLuN6kjF1gDGjY
+G0a+FT+agdEUkB9QpH/Y6rsswGJGnydlXc+hODlRPK1AbsX/1vouK2cDMvdlr/CioMc2skGxSCG
ldCcgByB+OMlANARGUkJqsb3lV5krdig7/vK/Z3aLn9VL111mXLG+5f9PT2lqB79a6323NQZbei1
3HLCHwbpV6SDXoD774mw8IE2/Q43S1Augopik1S5MQ5yFvStTT5JsQH6Gk7LgYlNqpEKRmCCWtPr
/dwVxDqHwxDLNC6HyHgDot+BpKQ+wwgTDEJfRZDSOTmxCRkmSjNeajUJKKrh1OAie55voigM+XVK
9LA3vqx4nrSIBRUCFwGQ6YqEa/233WjiwTRCIInndyvghH1mdDt95TPdWsEHg8thM40C2nwrGWa8
y6N4u+NOkFyx/cGVYyHcadq1BZeEfWwSAQJcR8IS0A+3MvO4d+vntfbaHVpKTxHlzztuXddn9Bk3
0xTNOuk+3VUaNKO4uRvlHQcXvJgvTIuZ0Wy2QrrQiMrYvFF55ZoEhgkJ4ytqfus0gT27B22d1QVO
1oCtd6NAoulrXTaM+Y75xnj4hJfmX41z02G3dMbcUrbxGFga3Qy36WsvkRIPSVyFKnyxEYdzAWmu
t9JTWHT+/bxGZDARgU9+Fl5ykcSuGGi+CYwLcHm/Xm21ZRTAjc3WJhGdd+2oKohzgSXRf98aU9nD
59HukIL1vxxXtGNbvAuEF+pmsv1LCZWCVt73ZGR1BS2/nH2o5sWn6ST30LNnRktqzQI01CADhMQE
/33PDufCyQ32F19EE84GwUysVPIKjk/h5WEYqxu7DGD9iTfaFBTN+EBMknOjU4my+fq597EUzdfo
D1ibi8O1jJrWx2JCkpka0iTRmzR6BHMdUSUafrn9UM27tyhoBxRHF+17EA8RXZke86H2HFuexb8s
rZ1ktJu7NtYIIl48WVdtfLfWJ9K9o04oTG45vTg28+MaVrx8UrjSRZUtkuVe9eD8+51yJTsvuSh8
eqMo4uReZwSNG18brX0vjkPIG9WV/SJzEBzQmbM/cRJhYs7YCu3ehzOdHgSFkngsfCDucLVFGtyE
lBlxdfYfr5KlHeb1kQBenjQ7iYgUDjaaV8UtRd0TJ/idEoEKpPCk1hPlP1+pM1PdgnaA/N+NSO0h
uId9T15jxHfsJDGgqTAWudPOTHyQQ4rYo2cVfpLN/cQ2irC4zRxmE/bDFRt/ImKrZqkyL9kMLfIv
ACKH5q3thDX2XMw48dKNv9VTyAeicT9Oqn+SWvMvrbM/gkkZPePjpOzDiRFG9mDyIMIRePXUVpcO
9OR2oBcWG4vcKUTO+4s4L8BgDeyS0rrR1VveJ8T8AzuIUczbqr0RdQpfZwDZdLjXIIKuruSpYOOm
W5+MHiOPPTDAZ0vqWskoYo5AauQb9LHm2OxZY5FtxOwDfEaFKiUtNkeNUwto+CvwxIAxJ/hdGq6n
FAiPYuJhtYiKcxxBlUP8h2arnkSX3t7BU0R3wpugUSTrsRtUI16UIxMPrlV5Fqg0Mi27T2YVjGag
uCz8uP1g4CTEIh2WvRvAeYvaG3GuaUikolWvuolA5VO2z8snb3RFbj7MjSASFfpnFfgpxCUX8cE+
dxpKkxP/6GmBE4URiSmjhDxA55f4PAG2Jsxk5WlmJ0UKD4FikgLRAIWkLUEAYUfD1hdW2TLnLSiE
DAhB3yq62qEXYvlizT840SiULU9wpM7mF4ksU0x5BTN0nKQWf24iBsyrlJtEvDbEtMvdFBdeJdfu
wpzxFSH4e0zBdwOHVJU46IwZn5Acj8sZQOlxWIsJ1TRVd08OZpzHrLG7bb1jrl/L8T7Cx60v+rw1
WB4ZtSvpa8KzwJEEJIIbS9yhHwXhgf63/MQcXJQ3gsHCNjYEi6MvRT62/HLdg470mQaNy/sD7WPL
JcrNt3mX8X8uqvb95g2EZo8PupEPIxJVmQ/KUIYHLHRI5/C1gPdPCZTrGAHzUTS7k+uxYesM/dRD
MEk4nkK21iSSWoHBo9w6nmgx3qehv72KgMS317XOTRqg90u1F39sk9sIwTZBWQ30Uh8h+UkDMi6N
Y2r5BJxgGERnQo0E8fFCTNwXIFfvvkR3s1vUcFcOsBFA27SoHF2A8hFQHaDjzxzj2EvLZKqSSxVd
g89m8jBpRUOZMeA/IiOwPa7bGRXBFm8+E5m9faqx3+/2gZoE2PdfbIa6oMnHF/9KonMRagcAsyLp
U78eLsx55W+TyJ7ISNRMfZhY4J3bnkFyRYqLm+32aF6rYQBiCEJzow7w4M3awUUcI2lqRX+p+/jK
0DZDRQ+CNH6dsZrxQnMkU/IDisqfO6WN5ZgEQt4VNNG+jm7L9ou3N+1zwqxYhLUFUVz+xQ6QJ84N
2l94UCs2x4vur5FSr2H6GAz1pY1DMLCnU70HT0O/E7PRyCevzJfSzsJr1v2P3gD0IV12QkKVT8UU
cUMc4GmP2Fq3cnEPMitUTyh3CvmKmLr+I/nC7hId+d4atzLW3CrVKskT9IfX5X1NrKZGNW1mQ+aO
yHL+iXk4o+bVqBudV2WB2QXUMuA5sdWPJDK6tssv6n9SD17zfQrs/VIHNVt3oMTvx6VqHoTXvFqC
uTkAOOmKc1VPz4gWrTXbA7+E7LKBtsvvP6YKWnzqp7qa85VKcAbIleuTo+SxEHWsFfrdfzmyuvWB
RlDN8BleDD20EySMa876gZJ8L9jRZzycLmotxMjWhxJ+J4r5Vz9JA0FvcxAfibJhvqF5kSHWYfLP
Lu4siwUC2Fp2J2a7ewhJT5hAc5h6WBs7ek3gIc9+hvNbbT4JfYtyqEa5VwmX8vNnMBDsp8fLkDSX
w5ilxLgBPvv5zCWCL0BydoS/ps6veUkoRUoKxdQduG0+zEzw+jZg1uExbpwPkTCOruL8CZh0deNS
71knjgFPFN3yti810Pw8b2CCDOUIzuSa1ZcD2dirJ4hypI1EUPDP8xENCLgP23po37urdwC/q83K
iZt0zKg+r0v0KAfrcknCds+f9MvoCo446AUQj1dQb6PbHTjJK11+tKWK1NJSN4uMvKakUse5WuTY
ITx9C7izOa1fL/IF69KjwnRjJ809pecb6ho6P1h6zGp/tDs8Up7UQNJdYp/0VOf0p3jJXKBN6pUl
gC/IGIPoZ4oC6nXYUAx3Yhvc7MAk6DtxZkIMgZpz6TYmtlhJbN8hRShORwGsDzMVF7AmXIUDeMqA
hHik4Uh3ZShUGJU2ql3DnJ++jA3BoTiGSEw7ASTmeW6oCsXsHdSRfVJ1gIpYL8iBwUspnGRPKDAg
xJ2bR/MgkMuUArCsqP+/pE8pSrLpXC7TMN/riuu2KZ0a44LvtrjUO0A1LARMKQdNqh9giACmxwXi
hzhCuy3zVtUpPxLak7Dsd9wmlhfKz9TVXtZYqNn0oyB/g++ENiii1rKXmu6/WUM2+ZPbadHEqDlC
gQdsBoxw/JisrusFZB9FTXBIou1tN8bcbfk2FD1fw5nYazNdPPhEDasNBnWxTz9hSsSf4eCvTV4X
W0ieOOZ6SJXeDniWQnTq9DN4S8EJczSWKgiSCIu09hNcUZmrFHdBWvhPeL4wJWKwMUMeb7bnigUH
nUJklSbkwZHu8IDAshXc/MjpY39PF7fI4qy+WkO0AR3EtUYWMY9aKR1vinBGVQJXBm+kj4rFeVDN
/i67ee4xqEqJuroJACFQVMujqtkDWrY8PX/8bvqlY58ifGVkLuKFOhBDxv9Cz3BcdDybtsOshKnv
v4oLT6nakdxdbb6+x6B1zmgWHjjt2V7T/zo1x2w5do80VYpEmsKG326ekm/wBbyYs0kN16mKchw3
ug+YqVvTrryvJgogDMN3Pr7hG1f/sAFNTTbHkFaNvEjB5Tx0TCDcQTLU9S38sjP4qkGkInHzFps4
K7BvSnXkzlHH5cxRGGS04Dd+p6asd6id/M/E1BiNT4Ku3lbjqlQ2AFgbPFOxVeYg+UfSluTTL3cT
90zGXbahIhjannNhh10prxq59IlPGARMdBYttzXmajeMKjbGjM5YmLTz5dJYl9kF2oNe4LjU4L1w
Xx0GZ/Do1hC06GH6JNBXrWm2P1omZ3D9H8nZ/qa/4u1yhYFNC7u4j3gri4itna3YAH5SMoox6rAc
ncznabQJ6zsgjC2JUeFNcT9VzRZ1nQOfEbzlC/yk3gZBNztGBI5CQcyaqfc52wKZYcF6VzVzgkso
anIngl8nn2mAURh5Xm7E23WOIHhc375PZJezcjov4K9WcExd3SKtXrC4B3ggEo1KXhFc0bYde69u
e0a+syrfuHiGA2zO3NNyz1SH5e1if8hrsRmw4J4vCmFqU4epqre2q83Fu/+HWIt49H5EGDDiaE/W
O6j22F5ovUQbZmfAJvqVixosf3CrPmumZeNQFW8yLWA2LeJIeELAe9gTtisrnB+VvTpFKAe79OOI
2GshQhgvoFNMLuKHk51CDPpqBkBaDtgehlEbZHxudvEQtRq5gpM3VnHBMTNI3q4TBMTDRxy3rsAY
jm+OKj8r6IONw9zcalxHj8Gny4q+IPjm/SlVMNmiZoQHFKPPnchsBBc/NUecaSfvm4U7IgeEZ5El
HSeDq1i8hmudXY9jxXrjWKQeOa+XLFsSyisq7bIwoaTpDFn9BPQ2P68rz9ei0l0DULvC3bb3vFLN
u9qoudbBN+diRdXc+dO3U4ZZhT+SnxscWPHQHgff8g+/gUAXuS4KxBAZbq6kVryW/jyjLYcdwlK8
Yr1Yyn4OSjN6WwWB00FG3WAMbBNoEpTDUqERgf+MSdWWVc1z9/WpFoJlLaHEE1fDQrGnf5EIpmlM
UKWFinVcKFKUPsRs/JH56+2IBtYbYL4hO6UMgd5tjZkb8HsrbGy5jVccsaFsn7lJgNMgF12GYLLB
0BW3j/ptteNQAjS81EYBPXL2jOsGI/0EZS/OQbTRs9eSvC2UA0RKvTAbsxO2njiIXHNNh/63+LyJ
2v/TaSBeuf7QlZhKuP9WleNo5z3dUK49mXAv0fngTp0SFchER058yFXlw7FiyQ+v5M07iS6PQrlr
RtlGWbpPRPNSvI5DC/0KJIMcAyG2P1JOyMaGQPug8LI5uEk4ZBW5JN+CnbHLozcNehPvLm2W/kMD
yFpRW3ciJvv2cPfYID2YB0ktU1lmvrbvG3bStMwjnUD2gqPAXcXdBU+qgbwIqF00ow5Zdz0vh8u+
mrJYTx6OQiqG+4fvDMyKiHvTXz9VpQMmpUOA6y0AbwkE1zu9O7yysBwHiO2GeC7e0iZ/lOW3Bnn1
Y8uwr5ckzi/UZeb//ybW674zt4DJl5TBVnc2oEFS26pBwRg0MBHGcKDsnJ6EcRTxNEVQRmYCf+kq
CODVqlz+duCyCCI71lXDd//RojkkQIHJ3vpTshL5hFWTp5D6wdTRBC311ZNRXoWoCv8YNv9J1M4x
inkHXBokquNAKOzJM1ya66j+bwCKh3FZPITe2SGiGMVTvjdR1fg6hWFPkhrTypsG+R4DgRGUoVL8
ZxSEe3Kat6p3AWq/L8k24geAjSchTHfBgCl22VvauPW2PIgskbZClDwdbP5EqPJpQbc8jTruVo6E
QDzR4mTFG0NOOymnmx2PsU+5VrghYUjIZ3bLcufzqo3F3mFqA01c+0N3F+H4dKeFF7Scj9P0fnov
kLjpQhicG4jcCbhVmoihbfuo5hNW6AL1uBoilgYu+9XrlrlNgQl9YY0X5RKnJi3E4jzWmbK9t/pb
JJnMSv3f1f6HnY9I64eUELOVGakkOjwdCUP7Zgf/ESnmyrNEu6WmNFgi2NktKa+mAKtJ5754/MUd
Jsw+NavUPuYF8b+iGOPKIOoZi9y96Mawff6bqdD06M6B1b8M/47JBoBdNm2Xqhb3Hrs8WGeMLI4F
WWbbDJIVGwGktoDIwOlBan6nD7HFSPzO75lW4i2Q2k33GpkjPKkG1J+S18k+pafsXYJ8V75IK8IL
xTctWQQPkQFva4mHhCfIHx7nIHDMaxFfzRbxdEoF6Lh26yGgDl6VWNDM29K+VBrTzCG2Dxd1hPpY
SMNvibOxwodYR9gbYF+qmEjImTNxbfMItkCSKgNVEo40HUxQU+e/DptoDn2UMpnv9+Dpj6Vn0WrZ
DkJ9vDauDeIk2zqE0PdTb0I3A0lskwSPE2F5GJHFsJJhQu1sIPP1fdzXBr8yIGBQU0v+0pnZwrm6
XAhfTspZ6QFBWnaldOaNEpG4cfIpQqwm+01vqKNQKBpoatZl4vCuZ1HT+/zgTFv/Rs8AyDAvSb3e
bjI2C8Mly0kfn9X5zEw9itIr3vs/JKSUDOsnYk6xsgbuEN8IgKa/JmSNOpafQXbrFV9kp5oTcrdA
1lgBYUbzjGOXvKqr5uyeSMoRXWMyY5ZuBtwC6dtkP+Y/BUR6BW40Ei03b4+jxtkT0lwSPtv7bCCp
X1UGgmmNT3QBlV+KgJe5mBJLVUtCp7qVv+AYuNFw+Yvni2mC5KGn7zSvC8n3/rN565SU21cEjMZs
JZg580w6T+3t/nAyfz2PxIKze+rmZ2dV/NcVxtcbpkufhhkEme4Z52JRDBXftFP4JEHOISR0E3vs
iLZbv5JOVoh5bGOXokXZqNTfe5/YjhKgpK+dWFPZ3lvkuL5G+BA6wzZQCFljKii+jyeZfTErhD0g
/PPPK36YfTaUTJAzfi/CN9Nvtgx6vdzKsU3YX6J/Tq8+aC0fgAZHaGa2P8cRhIDLO20Q3SQkygaq
J+3VujzbqUCk8QOoJUSG3WbzjIZMQcAVMZvpabhhE1LxhV5PFvHDQ12to0RcjMEKOWGrB/WdGnOd
uUsNKl4hJ/KLouvFMKNLLujcqTpr0bJCXLsNu7Su6wIroun33OjjvevTX7Td7meLPJVjjCSCAlh1
/VK0m42LNSLOZPVY7tQEjRsk3YZWynjpP63cxdpMYnST3RWXJB2ctS97EJjYI1QwX7h+c4ZIndIm
zqAd5OrkuBvr6O4TCdlaPioAD8TulLRUnnoMBjuV5e8kA1WVDKiqAqIsv0xFWWY7/5kf/hxftQlW
Chn0n7zqecGTNLDQL6seN0OiP8OaV27yvCqck19kb9AoVOrL9dag5Z2wHZOeaDQgjKsLQP9Gw03c
NTlZHI5D32VfK6XdpF3FR8rGGSqudnejd4niSyZFt6en46evwHh7hEb3qZ/YMIhg1a8nVs/LHoyz
//xDwzFriZVel/Zf2Wdg6Vh72Oelrgsz9duTg5JE6rXzjOyNG9zUa+6qFm12OwqWW4ttHtZVQAcF
qLyGJSdoSg41tn6SFGm1SYJ1WDPBrR05xjx7ndiYXsMnO9Wh7xEP/2bVAtuDAw91Bl5q9SlbZfv8
q1okop0FSDM2jGszQp1q7Nl1vbbrecYA/UtS5RjDWDNVfQjz3FYyo3kh9pFsBarlrsEtB9BHXz8a
Lb3qLHJ31iX+kCkLEg+S6EQeGByYglOeJMUUDmxG3Fwptls6aJ0qQpNMacQcZRgBZ7k32D5XIEs9
aH3sdqkEUOHCwUY5btAh3/rOMbf4EiCavIkcjXXdN0gA1PrSC3F+rfYUrstRBvyy0Rwz71IdvMuK
j5sdimSClkk6Cno2E4vA/UegCYZBAJwA9Lba9KPIBOtxFRg03V+Ip3AZzsztAcPtOdE8n1NFnS2s
Mk79IRDZkID8Athtcs45e1nUQ6/dZsEWjz1eemZnfVxM+wkpyho9HV7rpxPOwb2xE0rg+miGRG+y
cjwDQy7pOFYvG3mHhE32sY0KBzWgDhzEmxeaXqklNIHLDoVTbejfNz6mb6Hx7tEPm8dbcdct+m7k
HeeN9gw0iqtYpsRsc4W8B6QfWMnu/6Uy3Clhivy9nQDBizLnKE7o4jbkoy9obMfItCq+SIBvHncw
IN334juo6h07cfenRaZBDhMSUDpOusXS7QcnzozqvZZWWPgcJ9hVYHrnnh3VweLt6iyMzekoIyvJ
7kDMIp5OBfQJuKgFuFYRwj5AorAAIc3I1W7FJXe+1vZUZ6c1AJWKFIIqYK6FimOeObT1OzxcNKRP
jDpvNU8Y7wcF32EUBLx203fASjGRWqRaeXiCDTsE15YP9VB+O/yaG0BEJIG29H/G0IDWihRPgaMv
vTYCLT7o7yftfpyo3lrAIZD4CkW8SHqA9WpBpZ6VkOpy1fVYA65pQA+a6IDphoyMllgPmDiVQWnP
RXAfEGf63lRlMneLn1+29dYxB+MYsyoEokNw5zccTJteGbkuxoQArFsMfqfATcyIO367SlaEcgUC
wME3esR1hIzxQ4NoO6c3B0VTNAC8ZDfyrBaf2OGfhtCzqIrNgVT7SqJt27ZjZd4aGFboj0RsI02O
HntlxDbioW4+rWNv5kAQ9Zu0iKxXLMA9s+ykmvC/E0RBvUVzn7GLHjUXls+ZqAZHswb2rknrNr5p
yfQSZePC2/QmkyaY3EO6nFdAXks/LLGBoMwi4a/RmwQFrAYl0z1nFgUTOYxzgppcvbkplTTgu9aX
m9NZjwhwEL+YHWqmPyPI/hbGvjWel42SPEZ/4RQE19HBN9KbSlq1QGNpOBCYAI8FaojTPkqqGeKT
epMkRsP17m3e8cchbN4hIJbBCIZseWMZppqczH4mPUPiHD37tkWhdL9aJEN1ggzeYZB2t3C95k4O
xgmByf7n2/I3EJ77cOM12+UAIDPU2FIZe8BOamnah/uQiV9jVYQsQWwYiExOZgeruy9prnSvh2Z7
kxKnJBvBOLWDWrVPDQtRBlAu9ADq6RkjJOb3kp4QP8iZ+MN0qH/8CueV0wquEAaqyi1J85HNx8ng
kr8yGh0+JG714j1CrTHdQiMrXn1x8+fEViGa7zPtfhDic+uA9aQwdryvslQmr+RnjX3MD34L+GDo
1iNq+GKsHxlDNafDs5PoYlLumVsAazBv7B9HrzlMMez0HgD2ostmQ6wU5XXngX8tDw8MIjbFwwUm
WsY9SE0WVjmHNVOTgZcZWdD7Ai+D3LDz/SBLfXX6rlKX2toUuGjlIPslhXo/J15odg3+BHF98VQ9
snAct8uNmaq/F7k77LY4FtBRHmp+7XPwYUdnAZCDMmA5IiMVlXlTkZzF5V3PBHHLU8eW0klHzooE
Rvo4K/T8XcXjfAHr9L7SVvOHf6m8ZBiMycC2zG4zFrSaH2TXh9d/htTCXQm//B7YXyVttCd7g5Qk
HDlurl/bModKe1DeSDBbYjkEtEcdfGSqkgUJa+TI7WNERXFnEXXTZIDw7gr5aVKes92IBKR860we
QowbfxIVAZyH/idOANvZ/7jpR6aHp0L50jzp2cZ2MIB9p+T2zMYdxxiNLP1d3950BEfwlvk+sH9Y
dPKZwWp/zY0esogr7Gf86iT+TL5uyyZmfIjcn5DVV//RLR4KVYhmtwAngH9rJrnx5cS3goqwQFFB
zKHDT1gWTFaZM3/KGbbK+e/ETy+FGnQdj6LGCkqkQnE7sGGdEo/+Q09YLdGK0+8Hx21TBCSHPCYP
A5lbwkv9VadPAY/zv98AdXqBJQZYkX87IIIbDojKQvx7XJ/kBwRKdYCNttE8i/wYyahcml8BNtDR
auLrhGFdTL4htlrtni2fpRiLMbeVoE2VtEarZZTaQ788bkj13bWthayLdxIAIwVx/qxv5hWkdDqJ
s5/tCEDOq3tKuqhG94NNNrgNZpRiZX1K9SK+O/zbF25i7rekHF8YSyaVJ/rMBi5s+9KxYoNtCqJJ
kJsLFZtY286rYBlhflddg3mcGxTRQFR2/VOi+H0h3+lE186OLDNl/jjD3uAX8xFsaY7qBaEPPI3R
fYgdJVRd54xrzevW8j6mf4G+PPLtviPLAtoZ5WI0BGFoN4f+v1UV1M/rE+Q1EMVIdRT2/RCsOyIT
597T4agEY8SJJheU4vueOWatKyEkmPn+IfxTzjyiaoXtmNZCKcaNyk2a5zgPkQpraQiqx8QjWNhs
eB1zZtGPHVHNZX/+A2seN0olCTn3W5cQpHrDHGv8ix41zsyfKfBLLXBR6wym9lBtAMF2jEJ7E0PS
UMXN1Q5MyoCvigkrco3jbajqxxLkc1nI292vZrr0qDPLNk7i5o17ilyBJIjxXvgCq/YU7macBK/O
buAsrsmvj0KvflvMy17YBOjB7uUF66HPQ72/aJsZ+K2YEyTQo72xFpZpiaDHXuc4dHbBvM9LQ1AR
9CXlBiEjxZvvFHw1OkrttZInuKbgcPbOicZ9oIe90oIu/npLPj7OFx/q6P6456ZYisodgtkSrp1B
dSxCa4aJ3URKiWL3KDDG+7hCFL3UH+505FPXOM8WDmW1oYF9Dw2UatcLvpvV5rl7aJsr5yvEEAbV
U5WybihQJ/tPlxXfAtRfQnTSdbdr1pzkiQ7ddS8eB/MkNvUDFaBz4JQocinvymMp6+/z39U7D2SX
QrNBWvm5y7W82UrBxlmKkIarv1BN0Y/8gR5VTR1HTCDP560J3sii55amfY02IUJjMAFxSo4nqiqZ
NdhRYXqIxYzeNaDPfW25nlDlLFRV2pHwCKMqlp00yqnXyw3KEURV6tc+prp28TyVV6k5LCI3hbHS
eUMtgDKrLVm3SMbxeQ+Z8LF7I7XnWN3LD8uMooJgqBcguCLKaBG4+vo2HF6wxYZamIi7WPS7qilT
3hiN5XT9DZg3EarbtXcfPsUm4Ert8tTv/Zg4Pf8NqPOqvKtuwUPJy0FWmGpcyVmoE8F/Y+oIZOf3
CxoJDdtfOj3RF+4pDaFHp5ZUdiyBBjCX+SnexoV7JAq0Yq7kAenC7u/nbsiXsxvOoLAXoz7b44Tt
G8MUdXQjniubB7xhKFvW35/C5LXX8N3lM50kwduT+S9w7wMgND644gjuUpHQTzFf0hPAxdGKl30w
ThaC7DCBkReRzaDDgwvAzN36hSS3GWwv8A3e3xe17kK3ixkgUm7rR5KVMonQwCSEgDP2A8lbjDmn
1yOC7yn5mKObWxe78YxjDaWCIsfXgM2yNpMx0qUQgxAMxIQZeQpgEFD4JO0aUfpP8/ytc87Uj2W9
IXsbaskuBOA3jEKodxkvhK3l9O5YPY9xwS3NLe+u62zMk2t1e7IW0rI4W9PP7od/BlOO+UHHqzLY
OSTLPMeYwnr0fRgU7EYWlQowgbNrQyCs5wsrV5diRGLPNGEuaGKJrkkMxHNy3NwAlv4lGQR2lnCw
QJn0y5EJaKEpZFkL7Ravgl4nsU13/EhAVVn6IuZKqDZNHScuJfrP+ziMfGbszPzyCDvvlQEri/bN
EIE4UXrjFuQs5xtsgzf930D/MBCgxs7Pqnt0RKfuCu+zJIaC3tIB+2BfMzCCsvjoP5QT0oc5AlGi
S86ZUb4Nls0em9Ewyrt7pCbWYmgstYtFsKdm32TJl4JY5Xh6U/rGD6Jf2Pso0juSoc3MYURmPiI2
HFf/Btfoufgm321J1TOXvkhsD+NIoFtXGw0w7HDYQqJFDIwLBKnBGS48ARXdAmQQ+69rpyYVbtjV
UGVlwU7Z8wfRvDWPv3KYUAWGKRDl8vt3jx9nFHgE4eE9cs6GQ0c8oi7S+BL6OJOPobQCDJeYs9uj
Kufru5wYxDs4BWo7Xvz/BWAJiLgGiKyT7GB3MpZLD+rGMYartkwQu9wHaH3gRMdg92A6PsfJ8ovS
74M/Lnk0tXI0Re+zc8dX/KqdXAtbG6evEENrIdFlugszB+bnfmJLmyfC+PkVwrc3quMSSZ8MGB6O
7+xMQuQ7bCoXeJThhhbi/PdJ2BNbBlYzYKy73Fgg/FXaLJexU3RJSRbKq7uDCLJ18D5tb0PvnmuT
lRL+LLEmH2UT+qUj0nO2r4pxfibCR/iYgZHktN1vluIw6Fa9czAjmszwCD5g9g5vz7ixFFqZvhho
Eyu4sMHTQ7/Hu9r2K2vwc81LHxyPciA9064EcmQvPDC7n70RzLH9P8xS8/SSaq7unJRTSCoVRu1Y
ruW1jkCXTyJgH2Vecp7tfiekeXmhdVNvwSpXuwiDi2IAmHRSWgrGmJO920rG1Eqlg+vBb6tFew28
1S467R6Fnz5BpiEaKfLZ+p3xCoR6LnxunJ7Ybn32n9fqyj13d8GxfQI7vnke6jjYDLM9cSifGiWK
D3CO2EiEMIwwAEwNnw4lZug/Byh9I+U7X+Bnl+wYjDbviT9Un79mbtst7TmLIVNDjAh/yincXADy
YrkmBtXPfRo283l68kmPo72m6j02c2wM00jauFd8vVecBdLjnitapMZGToPuMeUTVFb9HPScfl2/
Y6BkCsjnCBTWR3L95XLsnhd/0MVf0oiiwBV9W6rkYydLoRq2Laq6pHqm+OaCb0av1D7m6yUcSEOp
eLkO0bwTWZpviO6qZr9j5Am0r06D13clNa89IgraJWTaXjS5+wLROm1judWhvr7PRlRDguYYksES
DeoKhdPqrCs7KBpXFML8YjPE81LHj8b2nEZpBDu3aG8Dbq4n7omZwlMO6XP3cnx/Vuy7bdpygIxX
5t861f2RGInWFO67EtD7GspKCz1m56Rnvzk8ZVfJMyaAJ/CL6mjCExsFpkaacpEJprTvUmBzLlQX
ox5YWyzzlveluGjgaB2KPIbxtI1X8riznmWQohOCz1BmQfd9VPUuzlw1+VX6r9vfunfv0KZZw319
JSW+vcB02o5zz1W7W6W1nk6ovuTYJeL9Y0FjJGdAIQqh2DQAbCPy91PQgy1v7V1AKDNUwX7pBNqM
4fgMD5EGNkWVb4GB685tt1KwADYC40d0H8KKA5A+O3me4c9YeB0TR42r9JgMT4xvDyMIEBY8KgXd
2DZebnPU9XqhldRg+VJO5Sy62SxXs/UTVA6TE4viEiWIOJGYBNI0Ahn3WvvLuGBQI0zcxJ9fJcuk
AXHH28uw/AwG0MaB+N/ZoauYfkfIcsGT/j+BxNeuoXWOTw+YMZWD81JM58VzzwD1aJ/uyOeBMHm4
kpXOpwkwVPCLhFcBaOYY66hc0SB1+RMf3BojgHzvV2GvRZ4DYvv/JYl3YeQt1Ht7SfZ9jNDgvMHZ
+q/H1koRoKTBK3uVlGduo42fiZCcYF/f1lY49BijylIVUMzZOZtUOa1MiGhAdQwicjKGbdlzbd3Q
1Jp62YKLzxpQG2bEcgMqUNY12uyNKlFxF53mCFCytD3OLtVbISXuQvvRzthHRG5oFbD88Uj2SGhN
926h81Q86PbVcR26r8k7jXN9h3r8g/0+ItfNuAj0NMNo6ndpwEQ443Cpv1UzW0vVIQgmMZi0TZnm
OlR0laUo+4duZbtwOVKrY6gZpbx44QxyL7pQdcE24gmn8HFYQmbYXDx0U19mVMPK1X+yu8bSrOEm
BAxcrYHUpXKZXGSNzYXm7ZucBCdNlbIYiAIPekWqPAmCJ0u7/KeMNnnvrjNNK6bLIFfgtK3DaLaV
zpvn+NSZQkZMEf96OVb2NWdDvoertFlBiWUxCz+3WFZMxElvJwJEpB0jEtR6M33o0RkK6N+AoKB0
bJQIZ0OEBNY8rLuVIOrWvW70FUMDDRtrC7lZNbiCv6vcKpEfL5FDjKSjVThMUzOPbm6/m666lKLZ
Tsh5CZ3Qai/MK1sSZ6UKBS4nE4MMsJ4lpy1cAChi03ZaLOGzZrPDp7RVSwfYYPW4/EWdNfmDWrfl
Op8xe1peNxLx2KFgt+nco3e9e82+E/LDTisMCXiD1eiUQDsz8ALe33EaKFvm+VBIyWgeP7Raoa1H
W9ZkeG11g12doKJnvPj3OoQe80Kq1rmQTdrpxIuKSD1LJYInaJuTlfa/6ANeLD8JUgBT9O/XmIWg
oS84ax1ryw/xYlp4YONvMXiM97+SB9KUhiinFBwgO+CYzSIHblfRhAcHFzVMsdQI1YYcQp6J8gIr
oH7jPfDYMiP2hsy9Z1wEnWUUUDWMjpP7vW8UbS98fu+odXwjQEQ7/jTRGhv+XHomXju2sWHoHGtY
zdH6tkzbu08CFn6D7rWzWwOEOztQkhppPnl+y6bt9Ke7i8SrQ6SAEZAOaWzPL/db6zcMpqA8wAVg
a4uHZXVmKWRnILWxK6ngxlx9LDpIiYpjbYyddM0BzeekJ8V1pbbkSJq7aTAqWOO7kdyaNbQyJRsR
dJzNUdHR4oipgTbqPsdH9GXeU8dZPw4gEj2jFu+LWZKSCe39zCXeu10NxGSYurUwAaGI5BcvRkAL
BlCLotyHGDcSs1HbL3NZMdkFvNQJ/rVBVSUKr+F/5n2bL09TPi64byhrSsQoR/Acm+6MM35cm47o
chTyLm1Y3tIBw0EtHk09K+S2d17rpDAo+6OHGErvHPxKvdOcsAL9zygs9J01hEqsYaM5g2Lc4jln
lXkHntuEYmbCMaE2Herv5JLxI05XWVUHcvZ482KtayKfq8qRsnDl7w/yBb3wYjcgCG5IBiM6EmEM
42UplXEDJnmT5TCuyyjrf2GGNASKz5N3cD956uJ5o9nenW+Grt2HOeHpshWG9NWDxzLl5BjC0DB6
rVmdEHEQZcjrbejH4nNv0U7cilaQvG5uPXyEJQlty05JNlOKZSEwIbVy/8r2WCvx+lfuXj5AQ5M4
dyGPxXoaWc5L33aU12khOaaunBJ11R/ZIMd4j7qytZwZ5L9cn7fD/Tkr6s04o492IYc8kz5YC6rh
/3OQteUx3kFZPNM515sqcijWgA68QTiRrPAfYbYbJ/D21SxvXozwCg3RItqHMPu9l0ZSvICwUNqP
xaOiuConzPilSFKwtosx5pv91UvqZBq6ACtjbUUmE5C+tEOZYvXLQisl1/8HnzI8jYttou5ukgm0
zjXcsCTslniZobKlHEu5RQmcKoktLzDIMkWYD+hhA8qKkfeAHS4A6a/vidAo3M008v9ABGGtvGBa
RtWV7fCJvibEPFKDHFDru49t1WapBlxyLELnB9ASn5js5ci3kA7MkaWYmko+Pp3AIDDQVFSqFA7N
tt0vNkifH5mFXx/jvi+H+VOqufVN97o7atwwtu7OuRfG02vOqdt/YwjkH/Kkz1zo+tFxIffBIOv6
TnMt6ynrt+QKwvWoY3duYuoJAjDoMWB7cd1Wc/+7W7t4/Szozyg99cAMsJRHYqlFRnleOzrj4pqR
MGVcBHsH/U/UDVndDoddlvC6R2ZmYDyKvJnceFRl8PpLqeSvgAUsgk7AvQSVVL00BPLtdyDHEWVb
PWpUtMYH3D4WeuVLiBoX1Kwr3+8aFcGlJE6id//7WF+3GVTaAp6sm8tWI6LCrsr8r4Jp9SLRYyfX
uOyBQ9CFEXQUEKK8Avf6TgwLo1DRjwUraaX2/waPz5t4cJrDB/fEEyvhku43PEcP93Q9+FX92zQZ
68D7EHVMMRZEePC2PLQgNiuUYDyWhgpqAiVhYV5C7QXmG2LjQsm8veDv6SzRk/vP1pVHLwY1/Dzv
4OjPsbjCmF3De6WMk9UKWPl9Ukaqhm15ICgir9iYCU9IteytGoR/hE7Ob0c3KKzfjU4W8eS0OlvU
WevEO4h/2XjPO9Gy5i9emtYap9wUs5866TK4Q/Rqh02Botvg2teOuGe+D3OZ6UXPvvSi5+mQ2mlB
eej1TE4XwjKWEucEbHgGwfvpk/Uh21LEG8iS0AcBO4EUTTkSOEbWvX76xug917xVnORQAEWe8TSA
huT92O1yeTAbIEOMU4W/BjUAPwq6Mm/zXcCUoXINLgnPIu+vd9jF9vv5gOb8PbHDS2k/RMpwr6qs
81vSpoajDRAXGrZq+lMVq6lkBux6mZ3iP8qTMCti2YxdiB7iHKPoHU3MMVrXtST+lQXooJPPAiog
czKrDCwagykENetxNIBwtjfN9r1mMz9GJBM/l5KG1BWuUJBR6CKqrO0gWQMs2Ss5ERncupDeGgox
mwBecHnuZx4QfQU7qDedapJ6rUHzmXikt+1WJhb/aaJvTRpRWw7f3JnH3iPnh6LM5HzUZNdWBIWh
LNJkVDuUctzLZ8cOQDdqU/F+FsFXPMGuc4UIDKFSqM5sJ/DQ2PItFbih+9m5PU8sMLDwKTpuXFGm
4HkTZJZXbNX5D9OXulqAkyBoqd58KM2HgSQohgxhoTy1qccNfn3Z+xkaJkR/ZYS3LSDscGL/+VHY
WzadDBaWt1YCC9I8AoU3Jy1Rp4+mTE6Zhlyc7PFsHXk47Kje/8s8JjTVGSnQab4w5jEN6hyh9dsS
JYsJFcP7vZLT0XBkfeBPUekXeYb7q/Rs1C+3MuH4InFdyqpIkqXe4e7fN/FzFzN067uaqbuKuyw4
DOYyiiYJxj3OipM2yhSzt9dWEN6qX/tIGHa4Dpbq3YB9Mn+L6PGEN7XP2szh/cByou6Kj4QaPrTr
qjto3lrdQ/zc+CwVn2ZlNMWHQ4Nt3p+Uh5DTlMKPoECy0HaIcTTGMpA9O9sfKO+AeWYKyShW215w
BVf+8kYuWml0Cz8ySDtLXwdM+MF/IfhWvd2peMd5JSj/ECJxX58l/FO134ODbyEtceKdld2mVF40
LJ2x2CzEUgjbRkht6UgQMo5AfgpxJtHuuUoBa//rwTzip5LOOPdS4NioOZtumWMVgO1wsV7pG2bR
jxd8y+mKcJUBr19v4RmnMlXkgr6/KbLl/yEX5prIG+BDqXOYNFk5tRh3V//Mfkf0SOM02RvlUgha
qw3jOb67/vWjcWciaGKsWIgqZKmvzjYWoD6TdWkSTCzkZFjbpC8lS8yNrZsmqNR7AA+Tulok/dLt
ZeildLczaYbNTbRNLccP0DQlRp11L7x54qHCHNCLbvPPSNvVbOtZJ2rw+yVjQzlOzLWDrC40+GMR
Xeh4taGijS/ZDZ950XWi09WJdRjzS++6sKDHZwLnrRyGHe5F3594S9K/5eYmIdaRQMXPE28CpC+X
eY2BSBFjqupz5Rg5zJG36EXJCGTU7bEKsx2C4Fayyu8PpIrYuq5dBqkqtTniSlBIBZd1a6/clX79
jeODUjiUH+6F/9tPysUebPkqGVLLmAl0Bgg6chz12ensyvPjpSgbGeSILEWftAJYCs4AzqS6WmW6
lAsKkNhUL7nbOHxWPnfIDM2/gbIVnNlGyN4n6Q3xDRMmigisngT56yxMK403udzyGGb1P6XFFpjA
C6kymt5j9FOYBCewLIfNx2J3nprvcJkXw8Vn7K6ejVCPrlY+if4srvbfYH+wVc+n4/i9gGieRh4g
zM5OHQaxdWffrfmcVrJ08xntdfFJiMRQMnl1YOfbHMqKIGPtpTNT1lGXb2vupMH7uZPosQt5GCWL
ibzwR6WWEb/hkQZrC24M1OgtDcY1y0B6GVBtJ32POQeU0gcoCZgLuqFZeDzRKl8e3OmYyvrJcovl
Z3v7gWUhfMBnVMiqVM7lnKoxsvB0TYPDZf5PvxSUj4lbQiqKXp4U3acvlBUEXdrmB/DuNYprIDgj
vEJ8Fwm1kLSm282ysg5T0PjUi81IRAL9Zx4p0p98ou4Frzxnl6ysAiVRwmnC+gxlwu3JUVjMXrXn
sA8XWnGW9f+JZXBrooTeFMRFqbMoiHGr8QF4c5qE7AOZnFleNNMZGWd8Jfel5Q2c/LpavSornCkF
W/TSmgMDbXo3YheAJb1uXSyTJhbUPMM+l6VcNoNp9GRRrTvInXMXVJPMvLp13gjmoVWNYTr6PUQc
sZMzLHhbDOeRkP6e8XUSj769t9ZYVfqAPfG8xLsUdOrGuNeigkmSGYc6Rwp2ssqzw2LH5wyrY7XG
/77fTSj09hIoPvQAbOcuaKWmvvFamSkA7VL/9sOLnBfE3CvxHMynjSi/tHBu8o+aBc33grSSutqu
8c77eVmAZC1pVwLB54eYHjmjOtsv7MA7/k2I31Zt5ZK5irtmsgSNREz+oeuDHcd3YGVOgTTSzQ3a
l9YIYxhHIIpPUaKcohwjiVFMHcwo7C99/AYIrVy1OBNGlobVzfCrIiclz2/7e5zloyWH+wbwRi1E
H2pYfq8CLycnXHklGwdHPPJNioWf1STiO0j7tOCNuw+AAwcDxruzFTZe6RLDIAwp7KSX/TClhdoz
xFzGE5QxUIlN5AgY3J+22GdWzsPPqNaolo5xIOTPRyKSUFPdWJrri8O5zxgX+P/HlnO0ZgyIVL2W
cjAwbJLqWIz2YQGo9ahnsDCwZf4r7copTBeSBz8y1LUTm/HMc25dwP2O5CBigKZYJXOCThHX4bBM
1fEUwtF6y+Tt6tdBFhw1r3JWQ+q+MKdJu8sdz94UD0FaI/rAF4PCH+n1OgyC5WYMnU5LYnUnonYL
V5g9NbQdoiZwUQ1o+sRrm1v5Lf4dSHnIrifjp/2P7sJvSdxsz3LCUjNh8cqffeQneTs3nSZj8VD0
2BaPOyYJwLk51Fp2GHvtVPy0oAMyY41UUagVKb42fjEl6kn0AYO6uBPmfVl0A4IcKJcSYRI3sRCE
m+UFYkNo9NpRMRYh+ODT8hTtRrS2zW66TfsGEnZu0lFW11Y9paUz0rZudmtjJSggnEDcrCXw7Lh9
34tRwojNAWoAxy+wcg58MKQT4QRM1nwDgxJbLYGXOImeerVarGBusqZnKyJQfO7NbtzfD+OJFsoM
K/n7fQMM84aCbakUu5Igk6YhjMatMT1oy8scTse9WWSOo5SLxD/opMmhfYbEbX+6aCWj4xW5hJ9m
pmY0GsewJ9Cy7BP7PieP2QuoOstE4VxSkbY0R3dO9WjE+p3s6p3Iq1yyctYcg/b5jRbYHJm64kzF
dgxSW+4fGnTfRvmgaAcgXU41XZLxesWR9+mzv47o0Z5PGGJzO0Swxc0iRAe9GxnLhyveEDgMAqw6
A7veIoZYbAcxdCS7yXzKRJR2lRceJeswSMxyyXBU0RnJhLRi1zKnBDOKPyoKAupGBe6a8LX9nev2
JJ3eVz5cDJeZCVfFR+hqlC/XZ/gWcxAA4OTqqr+z88Uwcc9drjj6g2+Vpub8Cu3P4hcB8hhpNTP5
2jyl5MNYNvXnrLEBifuJbaHxxvZctxsUcv2Stx+YHXAHmROSiI9VHLf+r2y7t6gwhOtZGpzaLb9m
QDFZhs1ZkObzRYEHCXyJ4VFb0s+6iDRhIeXf0FxHueQwNBsAPRIteuWU9GP5p5XA2y6eJmFVJfkX
Semn8ur/1OCVpmjEalZpJwOBksjAyHerufzuplGtXyRxhSAtlxqKZReYEQkLrxTgwfcS/4Bp4Iav
mr0064OAU0VG87QDA0JJfbzJyVyM/xVXhR4Qlt/Dvvp6kor98uB6DffrZ+B6owD0x7qXUBfbDVJR
oeTBQNIz+9WVsesMWKvDE3hRYgWedDd1/RmprwZWdJIkoAcy6vQRH8Go6DDy3q6ktmkfW0IOePpa
+8uV1z2lLV75vQ7zyJvnuPgiiG99CZIffJUr4AqEWWK7ZTPnjkfx8JANwTMPihhUTbXHA6NH77zM
3DThCxRDaDbcBcQQvY7viyVy9oGYLRPrCq/RIWKQVd+jwN9snS/lBNYSZODUCUiIShREfOZDs163
mDYapFzZgCaHno7rSQ9qQyTEBsb3EYKA+eTHnMSLiROOu1MMKOVi9eNBKUeiJ94B+qXSMKmH9jVV
xmesdcfLSj0KErFH4JCjVt9zDOnFiMkI51tR1w/kLtNlMLS4o8XYO2K3BTFE9B6D2gr1FjHfX4/u
HzoD8tiZVNFpo0wMg4QsKZs25lYryOXAgyu8igh5FmTyYgTOq1VAuP7SYnoXHyaBKZ/iqb15lnO2
QN+Ho16oYJWFpdnSzf+4EbHpmyRDiAF9hMfldJdyjhtGPFqPtKRnfV3hRlwNVxyfPjCcZQQs2Yt1
uiRchv8HPjCKgT4GGuYmSF85JAtNbKXFR955Phrb9gcFE9JOHTmZ+u1B4s9SvSmT6FM+6Vt/RKv9
0Nu1UhMnFxAjfdSKEK70cg9BuaXWpVuVjf2XyvGD2xdizuEr4ug2Liz7Pkc+AQhLmmSUdrHEjHGK
7aoSgCXVd9CYYz+r8DukxXYkwKzAlnr2Ic2SeC0gzZlsQ17OhMs1dFkYBPORi5rYU2nc29TqS/W3
aP+tPfTlI9E9e0OoFpiuSQN+Bxfkjv2i4zN5FcHHHPwcdT2WSi25JMaxLeWwzLyP8HmoU8/F4vhw
ZYuXCPzvVQ5JFjIj2/FC81pgo7EJgjscrQexweVYQlnfoFw5qKEJ0tsvpd8DbPWaKF9ZYL/LPlz6
d9gT9Gec/ZXrMeWMS6YIf/nJfy9NzNOxWDF/4WFJcyW4nw523okMU/aPbyM2qntMyXBgbn1T8Xyp
oJwzC4B/wBagPv0/3RyiEnYqfcucaGmo2eHP6oMYUI2Psi25VtsGmVSXGaBp1fp+OjnVz85RpRQD
bldIM1/lzE7AMbjSY8CnGpgLFq4PPW1YmPR3Rmwsihd4gPy8aoQpdk0WDH4mN97Pi+F4DYMXlhcx
kJ3qRyKza9h9hPbX9UpP1OnMFV3ZWCmYD6RUz47JN4/hrlpdEvIW+GCDuaEUiE6setP7L1Ovp2Jd
G89eaa+/sM2myCO1hmxs6r2NEVzFEcloZbUPlz3MhEY1erOE2c+LyOXzSFgJ6xpoifGqArGXyAwg
WqML6OlS0mmsOLjRQ1cnmGTCNn/NoUxZSRVI+l4tliI7+a54Fxqw3QTldOhrXj5cVmK+n529znDG
SyTiq1ycu4WAp3whrCQGMnauHykzNYNsm47AeUg2RLegST/YSWQdrRwXOGwl/oEis+iBiEBYWEXr
pUrL4ox9FwNafoZbKh73uhfncTxUbs7jU/68gn0NHl8dkGDQkzUGkaEdC/JJGMIo5+OZbOPjVRwb
SMQLi29PfQtlx33YsWqZATMNqqeAxmon5aefaEQUmb/LlSk4ykDyMEB8qJ0ZCSrgU9xXVPwrJnFn
ZdUP8a8683FU9UprIqtkrH4fKe1cIcCB++yfeDLOCe+ZkYVTdNBIcIeMwLejQHc7tTVIWd0qiXqs
NBdv9rdXgUy/c5LBkaQ9Ja70tmEm21Xn3AAkYfUlHIVcAzp7HwD88iiZ6d0miTE4N8H1SWyNhPkw
YkB0uJmPFhXodSdM3ScL+HJJjq4DTZdcI3xjqcYGro2osOiM0KqJNxUCNZSaAd0OWSvUejIRPTNf
RFYlZGGcgmcbM5dtijlINo0f7C1vMyhhDLdGrXcaWRnkFRTTjLgEpRIMxpdrlII1PXsvnRojeGA0
MI+weADiq8chj6eaUqlTib9/nzBniR1Luus6qA1kSsL3f2FVclckkacCNicjTgFJkzP5SvuPNDQ+
NWECDn8X/K8hKgXhk9nZdsRYcOqkx8FYmtVH/DGsHDb4EF7Rh9aZS+CGko+D+HFIdfX18+gDz4Ce
qMtw+P15xn45FzZ5qPgMt1ntJiwtVPTpRzWMy1fPTaWI9GkDiw2Llh0tPTOKauCis7nN8NNlJVDo
IxXBOusStyEOmLHDHrF8T1CgPeP3fMAS8jm7kU7DVvPCK39WZKCQFdYXvsvO7/GINtshjv3excUa
YvDstMg+IoNQ+jup3Y+9BVe4/L0pvx2RowkLttNJUzrTUi0LqWMOWV9mlztaz5fFpW1MEz/QsRAM
o2lMXsKfddhsDxJDTgaWwAtD/UE5bZjVL336Br3d3hXGCpAoX253ZIxfHA9ABPlPJ4K+TltZ+21b
m0l1pQJFTqwWHORt907sQK8BrFT+kNRizCrrtK5XxEqn/Z1EV5t/Oht+NcAit3Z6AigkrA0PBx8w
+KsM7NhSQFTYljOjozAwUzZX+V7QdWdix2ezP1p8r0LNe0OP7HLdOikrwS5mXKyr4msoNubXyX0x
ne3p42mIeM3hmeG2Lq0CNiWDElZz53SR0HYrd8zO6bMuAcmiDqgZ/49U/6uYsyg8dbyvYaXpn9qF
UprWDT1qBRiooPcpMsAYyWbBGL3odT6Z+N04Jc7I+gXdLDG3eQEqQSypIZ0l/6i7F+rcPAfBlfR3
uk1cSsYM7LEEpvkyunIndjU7kJOBGv2vMMOMHaL/FIcVb/AUOAQLHdp6ZlUyfgUiJ0gpL1IhTC5+
ndJBztceRLtGRb830pe1yZUu5UHjYCoSzCWkU3Brg4dMK1gG2zhx/0ZITbI6K30O113OomAc/VLn
L7Y6QuJeAOxsNVkUvNGo8ZLVx6EJfjktVzqdO0rtIkBZ2l0gjlPg1Ie6S1rZse01YHq+QQoSqBV7
C7gyyXtSzH+2G/btg4FUXke6mHRaB2Sxoj6gF6iTMorDCLTAhuTIq2cDYdbmoLkHlriGSrQKUAiI
u1p+gXsVpTEY5VLiSrdwDQ39pzNItydsntlPRsb3u33zUzTrd7TNmjKSSHpwWeIHamw7m2TwOS7t
TnA2fA2hByH9oK/TyGYtA/CbHO0EMBcRz7/9VJa7S7LAYxmsq/N3qYWPNvyuL7stb2jn5geVKxZr
pYTUjGCB607K9VaYKYK7wyC52ra7zlMqUj6+MxbiAxG50XQoAG7mZUPARJV9e3QkK8b3tR1YSVlv
Ut/dQXiS8CXOS1vcpZe4RUOc+CzIqwV/PRm/a1rjFChi8+svBknBBJ8YypO+ctcJ81rpIjDXcBYw
T2RbqJtCQT8Tw6oYzbBDPYaFQgHoWKXafWzzmXk6jh4RnQLnhwTo4c99c2ahhmiaKv1YN7AfzTCW
aimZCNy7hb85CKsp5scSuluj3FdUAnGUy0XB8RlQUrggJfGuFzMPGFD3n6e4sgTZpTzIyoCvEriw
1q8rDuC3hbeAD0TM+s0TP1WDwOj0VNDLELLu6twi3bYZnoujMwZYJy31jbbGMtDJZ0tQuATFuorv
mE9vwT+VlcIPG5f7GC4wU+rbBwfF7qpcJyDpzEMlac/LBgi1wLMVzldhu1Pd79R0tqIpOyWxJW56
OP8i1nU2JZkcVtr1Xk9iAcf2iT8LYVHNjprlkrCD5srfm34gpcJxOEQYKsXcnnqaffV5heE3OGcs
+tI6hecIFxRGOY2Yy2ULS4iB1EExkvR0/zeyM3HkVDq6SVTAGChae6VokWrReG0Jk3V+T5/64lkj
PAq0DXZgSe3sF1m5OJGqNGvlELqToj/WZ7HOto7/79zE6+zmtY5rOp2nQp36cz1cAf77pBJwzKPm
LTisAdkv8DD9ZuRH92BOgoEKkdYJkUYak1xl3jMSryy66shpMDzHyMCDF0VS6ATPL1LGSu//lGLm
uC/bEWVWy7WJ8cxjEMq8XY2DmgZe38fLzSOhhtdRt/rI9POMflBhPhoou1MBOe2AamagYueh6GpL
crLJXaI9Y9XC965GTDDBjrL0q7fxpjNE8hMqxLzMomrUDd1qBlbYo9/URdKjDrcwrbzI7mHqVZaI
XaaoepK7u4uK5sqmpcEhY/S3zAW37mnIbt/0YU/wxj834bZ7YNVvwYRNc5TIMlSUANavDhtrqi01
aDBheXUhNYEGIMxkAU2+q9msgAm6Ld+8uA6HWf4h5kxos8a7WEfPAn1qwWni/+9vUMd3nnCmJ4r3
R7B7gJUMDc4N6Om3hpQZruqD1ZAk504vlPyxkBWTl8vVp1ozPnRWln/dgKqTlm8ivvxRS9rGukZi
gwFKhnJ0ICHmkbUR7sayHjarfMJ0Mfw6X34D1Np11zPynoGb67NP8kS8C6tS3nM6VfrYjKTICkyv
fvko3MC/P3mXgL9VGF36ZG04gHtFmk8/nCMo5YLpMHKVhlu/OWEcv9j5TVxFKQM/AyxoYtqvvwUc
VePooL1MoGIKCB2vrOcPj8Lyry4zht3IyxGzARiN1iolWjqUpVAQLo/UF2+UClSUAbf9yhoL2eM7
6E8kXBdJJ1Nn+Ky6A9yl448nBHi1/7vxov2zEuH4Qx9PyfUcxGg15uYQeBZsazTh7EifyOLhoFc4
EvyFa0CFtuQBoriIheMHJLAvl5dX2zqCZsh0XLuA9reGneT0UACdJMrxRw9Y5Jb1kzdMQwBvsdOl
qd6ObcfQK9RDPK+a8MeVwcoZIreN7RK/8ufCbpcYDdiQ0gRfZoFKJ3vcCs45LbWd50Tu66eNX4AA
5aDp8FlT4+73YDXkngBSKxFRPl70zVLzRwVWzeA0D4QsUqLji5iRhsQbD+lPLleRlvW2/XyiOblk
gA8rWC21SyxO2ZZu1mDItyiEB0L5uBzRshacMjK+PRI1nXzD7mZTt/gPIeZiNBJXD8hRU1ZagcT8
kCYedltL2xcmnxFbNFuePFN12jVqVPLYa32sAX+ixm2elXFqhCNyg2USocdPP+jJblm0ljvPBFrG
qdeMlIYJZng7UprOTRLdHAtCLabA/4B4GPmmUQSuhaAWr4yjxaGcaKJC5eEAHKN3lhfuBdekew+A
zVkOZp4oSTztK0YoRFjbFM2KUNeyM5jfcweqE8HTLlT0Dmk5ZNc6L+5NDJTsaZKxJuWqw/vEpU4o
rQAnwxjS1Rpb/49ljSSxzSrMezkywj2OtrCqYLRp5BBMcuzfsATS4SJfuo27atalgZkDkroS3YNu
LBER6Vo9gotho36Vh40vSPXwQK3iQdZh7hR88ibJKgc14P0PbcnAnJzOUeHnqaLg7a21bo8+gyW2
joPX6o5pufdSaRFGTNm8lrroEsRsOii1OJqJUDZJPAkyScbhnIw8W/p2eI2/ndU5gvEb+qEvoHcO
crsKOgRLcQjFoHFzRyZ2m1UMcs4wW2DhpTOS9VLX3TPSC9XFDy2asGiJ8yNMuMQ1UnHMosNrcB5D
NnBrJ0OL0bzHAlNqvalAGzr8IzielPSuNreqvL6kLFqVNoQ/oEZK3LlR79V5GYKnyV0G9QPJzCIq
4IW3mUVAPmg3f1FHrha5zYvj6rLadeO9sL/jmzNGR/6ouuo9gXHRfV7DIaNc1rrczi9sU79HqYpC
83Icb94mDFJNI3MJvlT10yIGJa9LA4vRZQZ8PENTX6G70MFl016d7cAok7LOTvkOU699Ilo55nfb
UVEhl56DYqpENE6J0RQbB+ouxJWYgp/4FLXBhSocuVBwrVzO4/ryZ/fTvs6/W8+rS+40OrbAp0aP
gb4rIHCmfaIj/Bg27eFf33iqgY4MMKM5UQW0fi8Kivn75q/q0o1QeIsysOCrfT7al3doZxsrNpO2
Mh2jaliS4NAavkHuJmrzJIFnHWSdpBHieLmk9C3e6peQLqBPS1x3/uMrIdkbmIlmGGbjbqphdKnV
0NtK077xnNFdKXatQralzWT+9HZWebcOSIAxScG9aNc0UF7HRTsDJLpVmOt4lDw9bCCIxTRKelSH
Vgl75z7IW/9BoN6gmZQFwA6Wz+BB3nk1wjmU7W+CwtXWEZ8mi+NSXL0hd7bLSxzTOAf9VVRVFe3f
/9IeWb26VqG7Me04HVFdi/3x/U8Kaz5HFPyzS6COfjghX3bguMggfH6r3g8I4Z6TdUYZHPmtwY5C
lndF5sAGPeZQRy5rbK4lcGnpY+FE+dWzz5cuZmuFuNIwW0fx29dE3NzuQiEqqwz7av18fQo1U+7t
Zdxdnx42VElom5nzRgv66ZdURAolXlXdcDIlqAiYQVcDmdNoNxYFVEqN3xHrqXUPc7YPdPT6WO6R
yYgF5NZEukd5eof4z3XQg3QFksAJjlS7sS8rNO4UHOwmyVLh99wGFA6d4smWpldMQcEJQY8EJ2Oq
LHjfQOwY2kj4yg5YC9oAsdaI1IhAXEIxOsTvCqOM/9VioZTJckk/SWJ4nrnq1gPeXxkY+rJJ8kFW
e/yHcv4r/ZSQE+NkdftFnpsZCsK/fV/WvVzlq3LmgvfCZp1gW/YXeVmv07FyiKVIhK1paUqmdreu
fwmA/1PtcIQ/+N8N6wUHX9aCsq5Im7/2+3pB0fFNEltLp13BpIIv1bGwDlBlVbcqgzvCidA2nlLz
dGNtd4s47J3D4inaCYjhJStLIUSkq3WhR9DtCaMz/AxLAJAo717ByaGmcZlOTIvNgXuZpaWyeZ5C
G/PtWQafx25jTa+lSjVlxtb6tKo1dDyYUgIjxwOdz8QZmUS1TYNSrDQxlo37FuSjdFuvg52mvEnc
oYd3F0Cnd007uPcrhR6BjTeK7/edTwKkgENgf1UQ7lvWBsnXPHIHrVmqwk7xLD3sWYW9Sk9kqj50
f1jkOYvvErNt8/YNM0naZJIfRWX4K3LCcB6hvbvktm24uNNsjd3hMCFOp1RVYQb9kIHhSj6UrFux
eKcGTDYJ03sJonlvvwUkXq5a6HAkk+tNXonjipyau0Qx+34haz9DpJru1HyvRqDtJx6SO7ILBE6c
lvaCXwEoMK2/e6rxPVeyrbO6ZmzGjkg2pMT3idMaF78IOgIY/1cCROy7q6RRpzeflnLfgHBvNo4P
Y2RbWCma7m23OI8kkF7pKcchNAOSuSiUzFQAtXf5JNbowZ8m8fuYXl70/vzV/LHqJOIcSvfl8ZO/
ekQxEB5TpzOHDbiyA5trIdyatjEYzkF13BOiISc0yGouZVQXHUSeqOFGe4ebvhZ+LTqDbmb8I94L
ZU1CM8PjDZBeYPaKBZrCcvSeRUHx1TNv15+/J4OLPNq1beuW8qxSDduML+g6C0PKLfDH/97+7bNF
abzz2FOmEG21JKpJK+SZ0bYuAAz4W964+Ekq5XM3/lOgXwgQq5uZ+vb3u4+pF+qyrv0Q88CmAVRt
U/yCwvlxcqievxF/CtWd0SsdA/65w4uQvwNJWJbPePXRH06n5Hdw1VnwkjehKhe2b491zAIti1zK
mozygzHbriOjBDHVhH3+RV4YotpTKpT372GRf5Q0Mzw3lavZFYYKepxirXVQhenv19eiO/UZ3hTO
Xd/CN/xXsnd8rVQTKiWLC1WY/pCd1AVpcHo5KrO5zJOgvFzdtLT30MVtjpbmlwLZ7AbJF4vNH/lh
OF2U6TRB1Xn5CDgDhr1NcUlhYFjtB1SxPi35WSdf116c4galwEjL5LFD2nK6tf+ZsSHAvApve2Ct
8VJV5qRz4vL6HrQI7+bIlDp/eG28EhAlroCrXtFCzFKJcYU6i5Vcv13mylL3630kbrlYw4Klqm2U
01Vn2ZdDJJxK+yTE9zaEP6tetXpzwcXDb/U/yYhExg/17sKId7nKiEseXc9agKffsSEpO6ngQevd
tWWCIIHuIkxskE+6XQ5oNZ6ydmndeoXTPS10nBWE2XKuzk9FPrv1IbzrvFoyPhpKWAEVSVM5UM0f
Mc3Nbzw9R7kkI4ZRX0ZMuY+QUuhIWaQKhpPEj3dc7PMav1JtA/j3v+86KVvJrvXTs1zimaqT2j9T
MCs/1asl2anYUVwY4JTIjOwRNZQjA945VfzBF+JPN2TfZq2vi/FJyLbtXA/Pjrb3aMc7c3vuAOTP
AGAkn8rIx8iroYhhVvjyCtSSRbVMo+78Tb73mctADksu8L9GzCJYc8WDQC+Xar9/w9JORFoD+AnG
Z+PupmX/N/+p2Rr5N6fWHAsUYX8IQYmprZ5eqf3lYePxI5PBj/ittLzlbqdaIBx04E8B6UlzzRGs
F+XQlopScGGCpz5Lx8ELizXIWCAq538oc4kDkAXBjd5cUQ6CnHkGjy80XHzHH+fbkzypi/QEKiHq
AM5COAFkM492D/t4LPCPLuUGvoM+sBKi7+oXzFz0Wg2rKDXfIM9bXq/n/2BlyJEjMw+jozOUBzTS
wP8efNf4rS85uO/xBRjkoDNh0KNS7TG5Q7I9vKao7B1OILKYDXpNXIKBl3K9+GY2gopo9yunaW6P
HxmmalgF/ujBNJFRJekyHuRpPybopuvFzdIq2AMKg+wjYXO81OR3pQHAE1btCmk3gU6MvkLeRdlV
VGOvICgaVW7vH44ast0+FgE7Nh9/tw/7X240vz7nq7LUVFOTK2eUTqimmeuSVn3xO4FoRGanDcmw
GCDOVAV1WVZZ5CqnQcLbKb12VwqqEbLeYYOg5dkQBvZXGanlHkjkmqo3BI2lfkCxL9JrpcfgVwhy
Dta7DP8CoVHW4uwpRrojrhf1iWYpqSijPToCyGoR4gLJT6gUrs9+ebpVZ1rWrb4BiZmqEnhF15Lo
gK1oSkAC0v3Woa4RYziVAi2tOf+lk2uvf8GyElW6Si4sxykO5AGmU2RG/t4trxdTm0WupKZk37s6
GYPGN50f786rCrpfySDfUFBCMM6F5eYgt91gcby/sfSjK5qe63r7SqECPxZ6TBKpciNto/tUgDIJ
Z17uVqED5X7lFYzDSuEzpbKO7jby3izo/evzYmQBmA4e5IrFkltDmon34Mi0QfXTu7HAj1xWnGOg
NkOy/tQijHWVhRhxJsvaDDcjvJPsQKQPAUKxZPO3uVnKOSsCaVREUlsTJnurmmvi3rLL+CIcC7WX
qaGsf7u3PmnRUKdKrR+Nj3nd14FtKQUbbwpM+ygqLfe5q9XCIG/aGw70gwLpRak72dZRAHJMwEn4
8TmyRaj4aDhH1DP/jZAs/Mn1z47uDM6SeB3nM1SouTUAQQJgUgBWJ4ZBvFQxt9tK54ZfNsa7RL4y
9wHYgx4Rht8l5TVBfgjnRJcP+NXceaoLOgeOIwmoZYnuDN92TEWUoVnnaDoqNpcR7RJ+1c7cue/G
U/Ck68Ekc5ERYPyV8rIICs3Em+O8vQeaFYoVvKbOgQB8JXHTS34PC4MsSSkCreF8V+92rlG/znTD
0yiGyto98nlpSmzD+aWtOeHMmIBDOm9mbQyPuVUFujJsvjWbx/UimgNJbbg7SDg5gSvoIOBTPJrU
8ii+U/J/UvpnUUTImZtmSfr7fBQTZtyJptk+6YsDwFcVfBtu55COTPWgk2NqIFrvJZ1UZXaP+NJM
NCAOIWh01nGb1nC7Po3W0OSaxYCQgwW3ER/lt4vBN/QHw2l+MvoHaEMy0CBsOyZqziRTdJjsstwc
zImFXPvuJ56L+2NqROltF9K1LhjCu7ORlu6jR9O0CCoNWxhq8459eonlsMrkGfRscZROwFH/smgx
SlsRh+iNnkRj3UZ6ptDPzXuHwuGBBPkPy3BiKlWtAofMycZl8FO6OwpeNsaEEJ2WCI78YGxu7d2C
RM9WC7kD2lp2cuBLhmbKUSkoceytTGE7cOY5KOdLRw+VBykOkXFa93Cfq+Vv5N/EARfUG/92meM+
uY99R0l43F1OIpxLORs15n8RkPs92N5t+ReUjSuCSAoqlvgaXada1vbsBv96kDOh8rn/RUVS7sm2
jwbmvGD48E5mtnVm/m6EpllCpKTenx+Tga//7lu+s2Uph2iDsqUYaEhp6SHkNWPMY7TLsuQs1eYB
u+tg7KV+tDLVZFWkW1lYSa18AA9YZZtmEwTEL5Dw3Ny7Ci+yosAfBOacyfJDG7HGoaEotdZrDYAB
6nvc/A1sXRnkdMPRks+qFfU9FB7BCH3S331St1XWPjKbzSgkJIzCEUc0SZOJaWWmKAT5hN6qpIO8
00wPGc5+0q0ZQPdk4BUd5gN2vtwD+TOI152d3DWR6WR8RerFQpFK0cYnOD2X7i2RDiD1naQEwUnJ
n+5BEjkt/Y7iY1ZR8KobkaK+7FuejrTIQgu/gDLd/6hASwDEiS7uZHKRMEtRz0CqiCwubpeNz5Yh
bAwucYiSexpkMpqrc5NZCS2fBoGmExdAb7wkMpvAG54u/lNqns52mt2awJBoqiMZ5plAcwUAFqKf
QAZDf6lMGD+A/ljNOVCjYRjvxDHPkPnuEXx7SKqBl/IheYKC3wLZFi/noa4ToJx1ZEXGY6RKheu9
EevUg3uFX6B8oUVtL6BzWn7ShQjGMjOm/fKHHF2DfeEVfF7zAT4f+rhQsq/UOPYabVAwc8bbwJvh
ModP8A0PM9piWUQQ6yLwLGjdu8/vzVjGxdUTyNQr3rhsD3/UpsKzlkB46Vf+K+whzn6Gsp0XTZCq
ljZqnGDZ2QQ3mcG1SXWZguVtFsdtBBtsFs4sFtk002AN2JAYMDoL9RJEAbf1VeF6nC78omLvSxxR
VMha1xE0XGu4zI5P3t7JNk1veBgRah4TO7cnkWBV5Y84uohDcDeeNiGM3fD6zecmQ/rshjlaiPCO
HvQZ8xlojnO5Phegod/VqBs6G/h/gFc6X4dOHCrjAG3EDHb7dU3O+I8+H90j7styzoemNHalQ83R
Z9Wmmox0zuZW5mkNdenpxeG7+8BXoIB+YtNDOSQGFDsThIIVfZERQTK4ksbf1iv6UFA6wMKp0rmo
vCMNIYtpqvGHqDcmOdIcBOVAyIKZ4gpju5sPnW3FBlRSUfOFrMxzNZuBskm1+Dc0RUSZuiOlEn8L
ktdTkRFOG14MffP3oRf/suHONsvMRfHg2aFt+flg4FgC9EDfwrugVU+11+Da/4C//c31VVh58H8I
v686NgsxhEdZf0+SwZqKOMjxSwh6v5QnbR66MkpdrOloer7gvmLNof9+yQAcbeDJxSUyIkzz7Uxk
522hs1edclOYAV3+oZbHfQVzwNpZk1SXMr8r5w7sP5ASfxgNpTUf7SNoCy270q6zufdwfY4XMGs2
piM6GNwn+62m63r5wB6ic9z2HNThr1LSaSlUPWuWURbccULlh0NjEqWf1BFgyCIS3JeQglSWJN6w
tTjKn5+k6LeyciY1Yf1YHxasyXI34tAYRSiHxfewJp/USxEpu6VG4f3cYmlTQVsWzSBrxFtiJp30
8vjjTeJRXun3NdFNf8+hVW+untiZz5ug4dI4y7mQDhiOSRmj/alXKwbCuO30ZfIpllNAEMNDGWxP
XXrAwLFFMZmjPeZmsxcxwgeqwB28+bv4AVukZYhAjSCJ1D2yBYXcM44HzhGtw3NUkiKlSaDzz7Ru
VP9I6+LycowNJtfiynOiA2iMSCFCbKNoL3CxD6m/95KqUALIGAH27Evt+ea4bF7fQ2gcveEmx/YE
5DyGNrGTbz7rD3mnxvLDJ/4eTmV3D/WqZDaZhYBf0vhRlZt5486oqAr5AQ8m5ukkVbXpDzn3+g97
cNfbbeBwfKq19CJAbrZ+dzImjutLBF6fA6OZaawLHCdF8AXBtHz0j/s9ZKNRCLDosYC0UMaEVclM
5z+TFKAqj9unEJOBR6/NRSLx2iqZOl+A+L1Ro/08SG2bjFUdJHzoLfpfdtt2lBbITwBK6GHmxRFF
iAiaj/mF3w9YUTG06jBP6I6yyFoPfx1WhX1+xeI2BD/u+b+4TWJgfirbWmvOqiNsRPRPicpZ8mm8
1wkc/H0YpITib16i94svfrSwGBPYQnf5PQMBLiDwe0c341G2xH7h9KchUonx7gQVO/GIsO1eDfMY
oPB9tfKr9FL3qqa9/h7UkwEdayrpY34gCX4Ep2fClsgTA0FBl3RBL0w5l+rmSIAViTUKcLNt72Oh
376CmiHH/hiB/4CAPq7/W8uj7ojeTZA4COW/TzjjTnK6IJVz99vME67D/gKD1aeIAaf+Q7OUK5uH
jN3d7zzPz337hjLhF8GqJQF+nioDlilYrjHWQ1eaehdPKOIBB4My2OU75qZNifsErgArXzBvzqOS
3VJl7+2uXw3LTMWU8xm6UVI9QEyMSb8tUEPISANdNhaRT/VLLL3LCY0CqdG55HhQpxbMBQ0U8QLG
jnKc/8UgLLUrkFTWIk/ClCUOzVOUbyuYIG61zvc+jwC9O2XSmbfo7ttH1axRraX+7oXCIOyeu1WW
FSJDVyo8/sSLqeKR+wmrEM75+uX+qLgo3BnTfPJ3wCtc4eM3Hjnq5evVYMd4HDCX+HiVvH9mIS1M
kRb5H8MfE45ojrsBP2dE4rYu9pIqJT1zxZS3m0ZIfGMtat1hSMXaXSN7cSUuTZIl/6aTpPQp8Wg1
MkMEXrWiwQcFJJvN/3jLbTweMRAVws6d9qdX88UOxPkjHYeOHhU00pjR5fIGC3BIkdhvdZ3JO1Qp
HDGCv5aEIfpDP7liqazXjKvKZtsF7EqXzkk1lcFY91D1LrCqMTMyTsLI7OY1nNP/GFk4TFNlXelb
pJxfoHtY2YRYiqTFsMKMNZKJXPxwtTZV0Ms9+ANUuH6FMjtdIOAbYZxSvrtYV9j91twGnDF2PJOB
hkDZ4jqN+M/FmX+rhG2mZe6dCOBu+UDzbmo8Pr9XXUjFL9lAkyHymGXp0B2luOTg8JDie2eXXXmO
KNhmvyt99ndr0kwBKpcr8GYRw0UU737PsYuK5kv+O3ZIe4gZZv8qZIe+Qwgclg5AIFKh8HIOoBgf
jUbjZpW9VXo+KM692yoUsYV2iQCGQLWJOyr8v6JVAMOlpsO8+b6+PgwWmB+xnxgC6U3b7TZwvELn
PsaX5VxFYzSRrtHA4PeSRcnwI+f/5SVqMLgzXZrJG3iaW63I3rXR/hoZMTCLwsYwqRwZcprGcVMq
gy3wr016GKbwyzRgkJaH8HsZD0uAPZZHaIT9eOihn+VPWm03lw+qf5eCgzsnec3NS1smgJEj4Sha
6VdzAy67vrJC7DVnFnkneCmzCNm1RJbK4ga5HD3w8Hqt6M73AxoZuc/G1zNYqjUer0FSijifl1sG
Dhp/cyhuzTlZ54H4S9r7fCoCelCVmQQjGtja2USOJlm79nBorg8txv8PKAJbUVMTbl/8wAJ/pXl4
0GT5D1DzRhP43grv1owr/Pm4kXn3DE1YLnuUfwnXWyIkJ7i6+ZHoVUZtpRIAAKBgKpLsJ9bSZHb0
jqOVjl8bL4avOCPKjNhxi0mqgFvCfu5bxlRRvA6uDjhEIxC6RZQ7xAu3s3Mps5TjknPpYMDAYxIH
GrpaVu2p65zHVLmD3D1+NMCHFX2gfC+x6Vmqaltt/MvMHA8KMauOILe1CslvF7OYjmIQ1Q9Rg5nk
JF2eVMHlnzOfzZ1FFQ+xLf2DPfWIAJqMAUz8g2OMkTxrN0wFS21gn3U0WU3PMYcG4YNtZCY41YcN
I50mpShMbT9v73D0PIgRj6lx9dnELcxqtZd7C8LJ68FEt/8G+CNHySD6/tWU7r3YzYV9mznOWweU
A4xId+IT/VCTVHmiOHBovgimE8Liv4Sbtbqs26IgWfMT4FAxi/xHxsjYJcZzCEH/AQX03I7JLit/
BPPJGmzUtyd+vcgJ8WAID8FAuIwHcUEhsVIEU3SOmVSuHrn8/9avv/TgKYpDrCLp32KqX97eu5YL
JWpxM6/TD+LnzxcYxtDsX2NmSBbLOy4Rgg4CSOYyfZd2RgvKVoEm5ZMZeGf852uT/Mv5Z8XxNoCZ
+d4xqpRbq02Ho9qnD/D0jktEfpbWnqMFkro4EFivcAAJfiqwCWXOE84adCetGXYFTRdQx5hAzdFp
iumgdVabc9BI1K4oj1chJSVcR6BSg+OIic+F7CA2+fplbTZBXp2ZfawKxRy/sZWeZZMaT/3KoajE
QJ42UJEMF7C1CffoaVRi4CQbG0wGm5oIsy+CHudtyAthMsb6zqxOjQytQAxM4WCw2Rr0PW2yPegz
BXdwJYFzASHQ0zsE/OM5v8yag1YeD0hrii659jomR88hUVeO3v95p2pW7a2ywX2ylW5bI1RRMODF
RetQwA79IeEVXptXO5WJaAcUgajiMGMCorfUQniIswcdi98EbWiIyDIdHOicRgsNKFiojv905GOP
Y+xdZsYP0oE9yzJ1mElez6NDoH+oJgSfHCpv3eNZBj1BCPmwt/bBHHFgF/yuZvJyAyvXcMYSeOHV
ZRxoTryjfhG2S0cUu3qnOTl+R+Ort7ZPJ8VN1mVjdrxEkZf/sdelnp/w9+mUt1tHLjs5Whln6VBg
9fd6HtxWsGWlq/CLQtqKooZr+rcYfEAg3IpImV89HS+s1HxwPFbywJmrzL/yjOycHKPAahnFxyp8
j2PSb7kmYM61jK+pas2q1LdvWU3bSEbTPS5K/onBxNM87peOZcDEjUrBtU52yutrFoAyE1i7FAxF
bTBd8QGYL9DKFnaqNxJVjv35nhxH92JJGb64PjmRhoumTaOuJL7rudFPr/8q22IklAi+nZBMWOg8
kBWPS+7yprtb6q2LV+B3rJRSspzNbv2Aiqn9xDAxLXK2v71IKXBhVIKvSmO/tTxlLGwAx2Y6kuzq
eysqsqYpXkLFgQKxpfkcqJYbses70KSaPhnjfjj+FG2Asl2LiV5in2KrFd/SAOv5plQqmSIbGPDH
7n+ErtT93tm5w1NXtmTbAxz2bRBRGMwNiKkn753rqBuDCFfc0X9poV39nA37sizBNkHqIeYq7gG1
XsYZ2hX8I5Ly/EzeXNEINomdLvKVcPakyfBqoWXxr6gYHA5ecnA/yGPInpZ187vdS1Is3vnbabIc
gPOfjrLM6W/Q/s11JS3WIzLlfF1lFHBJe7rojS3NmejcQPtWJrghRXJ7zh9J6W8nJZffj3+M1Xsk
omZc46NLO2DJQm/p4WLE2oN7AhrCmfOSJ77ecaOw7c1re6VNsNRZh4uwKnzw7bB//phyAjT9EAFv
5Rd+FtAkVjgVXcseUUoGFgW5YBNcRLVgR1upna4x2gjmOjHsPughXh/on+HcaUVPjMYAFXMIL50v
VmNHfU5m8hPd3Flcw6TY9W0WP1yc7GEtUWk6cuEn9TUcAIHcujmhYAqbmqMQTDsqhrlzKDSJONKa
2i5KDFkQdq27h0iWZrFfF1SEmkyzG0DlkRrAARLuJHa5ehMdPCDwQPZsh8NxMIHsfwsmJySm0goK
v8yDu1AA2Ho2DijwqCcMaJSinKKCbvV68FN+Gn3lqOsqJ9W6HorrgbVpURsoI47hG7lD2Q3LiD4O
4upMmuODREj3wJJzOqtjwHlBZ+dOWcON4bDbzKwg8VTW1RkYbjitvoCzDaVpEUgSaQYJbIPLMDLw
muFv8oRVMScoQQCmm/ssNsy6lbc9n19CO7i/HqPU3BGToWc5/PKLwfIDam3YxOXe7pTHUG/MkofT
Syb3k4CQX5YNxacLj0WI/47HXrCz9CbDXtlwW6X6ocpYdQZJqGd4ufw54pOMJxXyYuXGz6mnb+O0
Ua0kHMYxll1O1CDhDD5ht67DYjdbcdgHESb5qX2AYSZPAX54Q0/n7FPPaqsnVCRAM2DFgybXgutd
eCFEgfEAIS+E5MvHTfJnb2R8+6QFvKVZYGaQzMb4N2UBKb1/frHXcjExB9Uu0VneXYKP+QlVEDHJ
FNyq1fFeIAT+TPEiAAaWFFd+gJK8saiJvIfbzzVghQ8zoAedVNaRXLtc3mM3ywg6PzkkRvGTGlCh
iVCJcBF2orXYo8rjGn/xrCvSOHOJMrbEHnlEQOIMddPbUAxQr154dD4duxRK91yh0r+ovpFejblq
/ZFyo+N31H8vTeTFDi3pcnGR7+5looIShqNvPIyFgashWVfiTFSkpJYM/t3lKyuhT8xmLDtDTwcU
fXmrcCFNb30KmcmQsGjLUlacaBZaceYptp91h6+Gqzx6UTPMfd7KwmiARCBFib+7E0y4w5DBXxUs
CMGUm/V0zr1b6KwHRSJ3TmsjWJdoVh0WqBzD2ev1Ax+dkUY92qf0kIOkSCXhydv3M0whGX0oZkPv
uwptYGr5Wh7npSvhTWdNTY/khxrOdWUJWWEKndA96h/ondrFagYusF3JZD4jZZzOmeKMSlX8aY4T
0vKhuln/BMi3DVLLY+wGKTyG1T2UeTM6eyqMozp5wP0Ld1G1xgRTCh0jTHRINnuvRA/qp8UEuORf
+lkkZqli1uM5eA2V8zPO6Z9uFlm9BzIaXZvglycs8WJVoRyDzXt4DGqh5iWvXpjfZ0gKFG3ZccNq
XRwfygi4nn7vW3JUcUzTudLucNDKLb47Jo1XqgYDsjVO3cbUrkKU1fhqd64oEetN17L2vRm+/nlX
GKdHIJCc3FHjs2JtmOA8qmGe3CFDQA+9l+JlKqn71Zpj+ie+/7yyXFE80QeNvd0kZV5OiDHGE/no
jwKQZAPKuxUhQQhPNsStZaePMxKf8oTlmeDS4h6VNj9Gf46Upf+ygMhN6I4PzCUuJjoA7J5zh4ox
OB/4FS5XUl7IMVdUTT4cV/a3scSOLYuy5NVIBzuRgqQGlW8i6By9rUrhRM4W/Ow+Rpe5AyVYEaVf
GlsJ7oAwoAKPqGzaCyi7zSdUtCQYX9ajcqlhj/EGgIN9BpBxrNRd1m96Pdj+nQSxxk1OHEQk7nAo
LLBeyvV/jX/DpKT3vB6JtSg6aSwqyIPTKgBgV6tc7UotngkyuvAEV8ptuh/BhhU4m2eL9nxYLw0Z
Mwk8SA6zyewYZ6+TxAOe26JU9h2+HDCrMTEH6hfgatB9qI/mZqEIjw6vPv7ewADIy9bIUSuKRizm
sh5qbmMF1Wf5SyJoJMZsGXnzCakZOs7tnwkfTu/2WzKevU9L4CywBMGeKw9uGOeLx29c5WKggfYq
zJ2ljKrG7GjscAPen9k4o/HaisZ/9cbTAh4+koKzN4GcsLqh1ojIQHti6+ZITGflKl/RVB4u/Hna
1kuo5TwqTMunrkXdl/8mgJGEUKCVd12rhbS+pKhYZA0Ifp6IdjwGaH2lCODL7hWotvKpiRGhoDoy
XJNEMaTIRRQOttyqW+Ao6G5WM0k9R2bNgufjtnbGYJ0phL57uIIDek8bfzhS3IE+eAXJwjgdOLnm
uD1dUayZGmZJkJt/OQv3XQf6EeSw3hZANOF/D2dk9hxtmcj2mFXS2tbUybEMQMAcJA27RlbPEo7L
10yRh9eW8QayXXNrSSwJRpyu5+U+aWWeQkIGfl1xUd1cpxqmHgca3smy0hwyGh2t8tAVtXe4Pq4+
93faI4h+tCgkhFLhktkf9kUktWF3O5hTmyRhslep/ncRC91RuRwk9eMAHI6y96UeqUUo06/RJ/4w
f1M78A+X4/BZPXrx1KdPWenbZPXqje6YeJa2Yl3t85h+Oq/tN6NskxOlezFjlrRA+THuOKweCk/G
OjCHtNU90ghcOTPsux65wPxwUX+c1Wbpzy65+l/O/XQ9oJ6zHCbZlHzDZf38ClIiblLfXw+kSYTh
wwAMa/KeTDUNzYtyHJr+KGqfkURltCK/hYO1RFpCyvcon8Pav2dzzZ6gOVwS+geOn9wo3LYNi0AV
V2LzrS8DZp8Lz4ir0zBLRO8lrGhNpZD/i/2ubup3jzFlniz8nBSsB2oZ9ifIK9DmcDXp+Km3RwfI
4urhXdezDFj+uSa24sZjfY1KgelvIFG1Sj7BN4iZsOMnKUs2uyxvg6PIyHbuXApOl1QIX5dPHikb
iSxbN61ilOOxilOa0nk+ZjtWR9XXVRwSew6xdCc2zehjssHFQOE1E+njRolVQbW8KkaGGJjpMTVN
20mz7b5DY2rqweBSdkBbUfxI8ZnaAh13PO2z1/VfUtSZSJucAXBhvgsfBe5QxUOfQVh1efVTZ1hy
tPKixAJbh4zPnrdtFNKiCCD0YbApHMzhJaAUBJFQtbolUflOB1dNeKtDn+9qOBog/KaBwJQQu2VL
cXSrxVZvCX6YDB8gWv0d9OS/0k8vFfYjQCvn2POvahuBqeIncVEyvRNd5nLc/p0aEjQ5lk7EmZBi
gLpO07fQWcETYihAQDrfujdrRKVufMekPV3L4Bu3VxZXuSDiPx3JS1JgZNHsR89ETfMKlVXznzhW
iP//h4KZEIWZ6J3Q+ZXWPU9Bt+duM/g+aQDqQsnDBXAMYSjjZ8sLhutGbFG9gze8kaODuJ4s1H1x
XARJMRWlCnVDBsTTM2UJfLp3l5Qshe80RYMB/EUy6Zo/gF4JeFtenOBc9M1oCf/hAANMhKnXvZMQ
5McegEdpL3OayZi47DP49x/Ky1+jGmG7Av1Lg2E/cJKpH3WUC77mduPDNf6BMkXprzjp7a9D4vt3
W3KKy7aJ8HVRw8bXGPLCCvw1DnTrMacI3dO80Bm046Lk8MJwqulgkQLCYpqUzs6Xi2qPVxwGC1pT
EZCEuRqWUuadh5m2qegXhjjjuhS82wxlPx+fI5FhZQ0XEVHNBoZttHXF2d52adfnm+g6FVmsZk6S
ZNRFkoNFYDiHM/h2vfgiO+Pe6O9L9DROURbdRsH9Qh4fJS9fUyiNAP3SUOEnmUb9rl5vgkFNYpcn
gqaBV9Dg4/qX7hGduiLY0wEMWZor7OOFFHKbD3eIVXY5ZOhrjwAwRcWvIzN++mv1Idcak6fZfo2w
Bs6qo1OJit/9BD4peaaQAS7/sV2wp5y1dAxkvcekjH8Q7qJOWsq7Y6HEiF2kdLqKJx9ER5SxYm+C
Ek3Zyd6HlNblEqBUgwCoCYEEcYb7mcaKOG/N8xTyw2yiEZXvv76YlfqWWFGhwDsNIfc1U/DYk/fo
Pv2gpgawJMXLlbC4PYdacdCUDtp3Gp9OKR+cxbInSM3oYoxpIwSTEMSl2ooAc8RxPThYi14AbeKk
gxuSYWHiBblMcGOEO1pgOzRd08Wqw4s9ZKuPN3g5hHiBtKlj1ehqlpX/9yxqvn3HicySXQPrHz++
EIL4UckeW3Bta3msIEHYtBuboH8Cq6I2T45dOjR4gW48lgL2/GRd2XgimFs6tIIAY+GgGGw97IRS
rld3oE/gpYpAwJIZD6VockAZd/ajOprA2UiLEVNPBKkUPduTqAZ99RsFZj4iku1DsGDzzxrKh+El
T8Hzo8/5mddslaCua+cE+AcE+bWMgE4JsjW9Gg0EcpAMrWqJ2YbkZaF9tlNXTtKLr9xnv11h+N8Q
Rk3SYOgLlM9ADtqDrEpSndSZlk/vwuRNryCrQiKGS6WKOeMbg7SrMHsBE5Rt698C5lCsVI6gZkw9
kjZ1Bw3wXwgjZeeKTe2VvRAOseytv8w7M1jcKP0pTXtY5QMvV39A+mV6IlBZiatjAY40j5dc7Pyz
hwgMSJB/NN60OxLzPByy6JTXz1ukT4IDLV88UXO1WlgWfL8hvo+63wZOIh7S1R/8dPWeWxumgQF7
OfIEsBZJZpfz15EkqjLwEwfdgDDy+39xpnCYOdrznHRRJfbj1qQkIIdcLIt/HHQGbN7xkb43Kfc7
J2abM+6bkfLniTIYl7pxjaiiYA15LpFWHNkftSgVYAhFaBX1OapNNaTi1WsGYT18P5YynYCasOUw
iYtswdqjJysIuLSRRzvnyHFVoTD5tvHG8MGZ3rks9dIv0Yhp+CWorr8F+qz/LtgD8wpLgvoEfRp4
5nhk21XlDMqaJ7EXXNRXWmHgajuOhWO6FLDI+/7Z2w23oo7sw3uTalShedaC+wfjmiNibXOtLnq1
MSzJiIQY3QIObSw4nYr2CQG4vIxi/Fb3fIopgrUGJi8v/EpIhJOoz/sjZrthgkWYZQfNp4yMzGjd
F8r+ciaJeTDYX4h+LOM4RWyfJZ3pr1Yku7rjTOsIzDevv4S0U12vzHVsNpnMo5T1aFwIhSB3q8Vn
no2LQUmDT7nlGLkCSVbDyaWXXJs/B1PPYHipXgH1I922cuL6R6Cg6qB+Ncp+B4UV9CcoEUfOilhj
FFUEBp/UJ51FD0Ct0KhqEdDC9nHsHN2UN4zOt55+USldoUcBtiNMDg42FWdTcXQ0YmxM/3K0gfYr
8XlVucYeo+91ZXoHBbWoLvpvGEjRE1X/sZGoKgj0L8Z+ASAniWZDQEsJLOEgZpIrcmlxiu1NzJWn
d5OLOsDcL2d4bnGCoThI/5ud1k2q7Upz05TWWYnmRrf6ut+iFXRljyzlB/vTIo/Gu1avIJFb37Js
dPH3ftL5ALFMMJR/3/gYWZDKuPv2s77JFbkg0nwKzjd8WXY2rU/hkgy1Bzrtbk5hCqqsJpFAHTeK
jiEODCrnlvubtxjgZHcwTY4V4PY0Z8kH9UgBKUEa7MzHl7RK1+kRF5UafDoLb64ZhDqRbzjKlVIT
J/6BDsAPE5WdYmHVWWJuFwKuKuT3eWVJlgE+kMRwchKEF/+89k6pjPLy0TPuSQqLaR92R/2rUxIo
VokU5VE3GGyQYqO70nitz2khC1lo7skp/z/OWC3cbX6+gv1Kw0q98PsovnzSw/0BlGrK7nvHbDbv
5/3VgDJkie46LkoH/4CIK/TiY2WT9gqqoA98lMXF2IIAGPoUq0BQi7cal/pLSMbg1gilvdL2xUG1
0DgVpe3y/aXCK3XcRFcXBZHJcwbibmB7SWS2qjCgrf2nVzDvCAhwlElHrMWRK0hjZYb16tdfc8xa
doVEgHwcNzSkUbBIgqIf57DZk4LqU4+lEgT+Aqi7ZK0x2iJ0tCh5yiLfTbKr0C4iyxGqVeFJphCa
xgBjv2qQryoD6mRALcaWPdvo781k7QnQyeD32s0smzOJD799gcjCCwsrycWqB989iNaEqDfMpz4k
PKytfoq24KXuicxGY/OeCYOlG+nKWd4M1ZQ++mzYz9N6VAR31Gzq9Co/Qo5YdgDQf5uETzjaXgEg
bsiKGt6LghRAOSzhEdMd6bJPQsquASuR1yRy7xlI9Ttl4MYnRItNphMEUAFM+tKAkdDa/PaOeAxE
pwa7ny3n2DGbL3NPOKBneDR2GVhDtF6tb15psp8vgvtsISeMQanB1uDZvWcjl2MHwcxT2N/bSpmm
gy3q2wTnpqTzaAXYK3EhR/xxCRn6tzQaMMl8J3jxEycWkGAacj+7+eZhMjwXp1HlhhtqDjMGZ+8J
S2zRmnGvQeTkIf2WIwqr7x8BS6BlJgO/aOfGrtrG9hiYWXfykp9GrOs2c70FHm98SEFejhZNFF5o
PeWHP6gqYT5Xnd1CRYIO+NgLvckJS8TQR6my/4m9PGMB1n4xcKqi03r+gEmZnlxZEHR/hU9QpgFJ
IZ52XE6umoYMseX4/f7RIrJknEyGLp90SjugfTaGMnl3wzFfRUrt3CKRG11f3fbAqpKquYqSdqlg
n+W3AoVxP+JOjYgudIQdH75nFD+ViS+TwLenMLHPMoRigzGoaGIfG6+De31y52SIZB99Jkd47Iw2
EHVoM+fFtGPWuf/nMjtUo3XYtTInhH+SH0nhGEhmYYMssDZOZZ3elbiTOisIu7miydPz9hNjoNaK
QF716hS3pVx+hddyUh2/84mabGPFa5WtIjsd6/hJ6sXuBIAtfnemvnY1UxhukywpY9W8/zZIL2kr
xkpQKwtyB96UtAPDa4Lw9As9i/nIBR+qhrP0ymPVFZSPgOzBlo/BRimqdweHzIYGBdjZiGiq6ORH
gKglYISCRzCDjwYZHBm0Taq+xJTiya8imJxaaVpprnqOT1uOwQoDpmAGHIugFCSbCAtODjIpD6gn
d6YzIU2sw0m9vIoo2HxQ0mWTligZGI2V2p2i2vWR3WQpAt0Tb7rV2jnnQb528RF5Li/2sJSIrtCO
VqFOiPKyXvwa2myI3pvao4jIfChSDSvupTKu3UT1pVkq2C8sd40ryBGbwqiFYD5jfdlE3IMX+dWO
GrWAQEX8L0Y43T1bBt6sXrw6RLx2wyYRTMZcRLU63N0anMEplnL/YGx5T/7Ro+43jIE2hW9hO0Rb
haR5xDSlWMmTQfxftD91Dz4JOb+yu3dZgxmWpn5a1+lQv+Q1NhZ1ZHHuGlGOxyE02oq4ztpM7mpB
Glx9RDTpZgpSihZch3zVuTTFdaHpGQrG4DM+L9yOuYiBPAWRjctMLlQR2w14K7hjuDx3WrW70A5k
4pT93Lyr99qNfRN5qpjJptWjGQgQHd4Hakr9pcnaSoGjEtMwmxUfKtDnYsNQb6SksqfxBviCEGLm
H7bHjeZ6zpUUyhx4+PdoDRUCUBSIDCrGa8L3tl2bVthAzqFZEH2qXI6xCNO66D75ULQkoaHaQbDn
GNHCh9+KsZntiIPyOCM/sfXY0y4K66bZK310MFQBw6FyN6U4Ryag9eLF1NEwqgSTpAvM9SdEmuyJ
Ct1X+fuZB7sRZwTIZLYIx5/kBJSPg1yEvgslP5LAv1PMm93HheQS5glh1f4rk5ks1cl2FZpHy1lU
mJ0IC7YXFld+nI8yU+osm9VgcU4xVCiGI/ItZs7+P2FCQAC8y7S+byHrxhoO0UJCPNGxSp6XQ43i
o0yvcW9mxNX6GMrLwGY/LzgJ1U02amhUICxyRcS15ZRP9KW39tb0xUtYow531sE7P/YS7yJ554Kg
KZlvgTb2rpLx53L06FXodkq69HEFghBXo3SexUivXGmzfFYSQWrgXsNL9eLFN0WI8LK+qpR0Ffg+
sgqcBy8ccDD5xkqgYkEMX8ZLNXgOjn2FqBrtGtSog0gHnUGheZhkkFTizAGM+k2QCSZJGzo3pBBH
rkoKBK2qU2wJXAnBHWdb+CKp396bNWu5vRJAabhbsHGWTwHABD2rzgTZW8/FLtnrHQWk2uQvyHoA
CW5VRR7fx9lg3LizubsbHkKEvoFJCqzpqNHs4KLdws/LoxCgVSR6IHQl3gRcuhmk5noMNqSPh8mt
pxu6HaIndWAP/fZVaHkZR/kaox4pMEIHp5hbyR4Nijv3TzZiF+7xo+SH7sJwZTGMAqIx7MLWqJR2
9SdlYZPEcrDKPOtTT2CWnRw1TE51AtGnapVUddYLJO8Fb0O9dY2dfxq4kzT5fRcxrsYhwxaMTlEn
BcjRgAC//e1C/tdqYzFTcbhMc4jJ03Id6rhCFAHjPB/rtn1MEVDkKIa1R7dPUK83Eb45muDA4hjv
tDVnGPKCW9AZTjaBI3cjB7fv3TNPQMZ2y5V0zhIcsBc/YbVTKzd3q2o+erxs8FAhMLlcDnoB+3DR
D8NJPghPJpt4vOc63C3Pa5xcZcYRNRGPErQberv5BmbI5IYXr/RcMzsBKIPqEujy8jDla794dIzp
xwiEY++9TYu3VXOHCdM5+kF3K6lY9MxRyhdNu4SlDdjd9tR5Xq+S/9B+gGLNWMyWMp62i7ClZfeH
EKZ+itos4BBvbcMWlWsMzNvr2xlLDqIbrbuFrI+90Wu58whHnbpSerfUQJNGDpK5CHaEDuTjmABH
j6m9m6ChfN7N96PKOgV60Gddgidiqjm5n5X7bTZw3zBNev704SCRfZMX9JpUwnZRseIB+8OrgsiP
CFuksJYU0JHW0CgtoJO2BBaFo2Ziz8G9dcgKO40lVsAxZ3aVwWc0IDBFpdOWuK+M1WuXiRXbaY4z
2qkC+KrnldKcdoVMUizUMAWmPkckuSx+MVt29QCHADGeP2yHt9yFAnr7lVW9JG4NTGgc97HJ+64P
SpxlEZd0ctOB+qkj6Oj3NDQ8cpePBHvCss0U0hN5fLGvKrS/JqphGjeSyKhXTrm0mGF4JiHzyfto
0qYsF9WbnDskb5Ipm2SXDEIEResxpekXagboYG583qYf54X+SRT1qvbExET6oNhFKnTsVwCBYqCE
nNgLoGEgywNxcFv5c1hOdqi1JPigM7vvLU25nYGw3j4DBLSwvs9YO/t2q+cznxDEA/Pa6mAp9oln
9xcDWfsF+n2QXfZcJ7vGVfoFKVY/yZPCxs/18HDwviX41lSM44Te7rXBu8w+WMeZnWL/qRgMY65t
kesSvECuD5roawDJro/mRNmF0gpm3Dh7yGQl3LbUsS8KS4/4qXmBXTSVSSATsJGr3Mv3by/rvZ5/
YbWvEWjx8owJaGq8zP1m2a3ABwz36ATFYFQXcQgfJG6LsGxF+rA5nRmdH+0wpJQgl20OenGz8w0P
QJxjqxq3C8Y/z914qkNrd8JsFQMJTQyC19yGMuf4wM2TTCOAES+KgKy/9w0Ce/zd4uzO32CVcQVA
3ZG05XYNW4em+0YOK3EIQircO9gMfOKJKnz8RjZ1F5nznVx9C6lgK1j8cQ2Gkhj+i4Z2Vw1LGycA
AleeOiY4vDRKhJVrp1FCNvcyzlKD3TP3XApi8+eVCMQ6EbZ8sYz3ia8dmXqYsue/63Aj3+Xvx2dn
vGHlTgdTiWImMNnyB/IVbCibrRVDh3VbL0rhYM5w3ekAVqBqxX2beNkgWpZr/xLIQMrh/QZYGEhL
uwTkpL72aTfVdwGKkN15hUG8MbmNw7xo6ilUnYpaFJyVYXtuRPEXzYFiSAeN3uIC9vy+vw8AxETE
eTny2DD1nmuAgW8HyKGuErsO33pbTu+TDYj1iUUuiQFMrKLYAMUJwzc1MEgLF+ZOgwj4pGKhDdrj
2JsM7Noi5PubBWyazdqRVrsUYGoGOAkJiU4e7S57R3iach8v5b0sO9ldZjX6q8+l/u+IiQjzMZxO
DCXkZUodH0Ad2lUIxwWmMc/tSx6ENwMUBr7GtkF6xDXvd/VMF4fdXJt1D9uMZmOfLzZCBC/fyzNU
cSYyH/kMrJBbAYJnQmuO/cu3fGgxpZqXE5tNo1YTYEjF0H588oZpctIg/nEQltAY0G9dSQFbKGIb
iNKLDALEb3Lfy3clSgk54bNm+Z2AoOpLe7/1+T6P7AtQQeysqm77jf+7/S9h9F6e+V3KDuEc9Kb8
dbdeJR9t9Et+31+2a1AG7dIKvozOmDeiB+UssuWMssl2WLWLJzJ4jiF7YDnVrFW6wiiHcKTY3Qeo
jMhItFawDWtZMVIJBMzO8m2rJJNBXXktjLeSjdv47f3Y4djHuG0a81xbzl9gCYfIl5Mgepm9qNV/
ms2NiNDGogo1PccUM3ZJHQ8Bjz4A4OLdYhjPjkra+0GdAX9nfQwxA6aExlZtqLnI53klTOXvMs2f
eTph2fVie6ezEa312JoL6MFz07WW40+6alUrknTejoywhvrp8CKTm+Lw3OHZH/ruE7Qj6zn5MK+B
ZCPmz8L337BUb+VXZMGOwZ5QaUwEVxtZzV+4pQXSyEcWWMRzCv56QCMk6CddL9uxbXeIPOGDiA9t
4eK/bors1tZ+RZtczP2XrKZpyjgwmC4Uk7IG2ueyuz6xCtiWyo5mLGZMuHVS4QYJvPAUXjr3xohI
f2jj/GdWVa22kWjuYd1INHYh36ZgfRJfKndM0nWAFbOv7AnjyaqvvnZwKnGe2JIW1zdmA0aTo9dH
BbzjWI/qz49txoiF1rh7dONmD6sMd7opWUPm/CJuxffqGCwbGepwXXYfuL8lYg6fdlXhA02YxHyl
U7SYJ87bl+ndjtzmIX0+F+3g5xZOiiiUugVmQBnnQVy4fXhxH8QkmPGT4aTlYw3jQBqQdB2Xi0oG
x2fGMm6Unjo0PD0MLKDvD1JyH6NqgsIOHgO9HeewLwPxnNNNSqQflXpdN6tM7/oapzewvX0T5Dcu
ssQbwdp2+/VluGw8tAK1ccvnc6tp8LpR/KZ5HWPSCXfnwZQ7lndjyBQKABbfKORBwXT8PUo/qwle
Vpn3v+xwJWPwTgQhpkQNPFK8ltagQf2Zc4XscoOARx5nBSy/He1UUFZvdkUA+pSOP4G1kXr5w7qC
/kvkirzzdyn23R3qiPx5RLEdGyZTXe6GqcooEWafbpQ1RbrOPCoEAv3avToctXZsGAzDH3VrMfDU
vA7/7uEWwNQyBCOwxIaC/xsho1noCGU44hDGdRVS5qkAdbEGTV6cqHtyaI/A0OB/FCKgiTzplnu+
M+X59L/Ob3DilvvHUcU+GnzQOLOhOEK3nXO9CvuYBw7MlMzwtEgEvGappPdlCuLcK75uTtXDdR9U
alu7+HByN6KXT/nUBvMDvt4np+Pf1sLSn48xTiTsfdbhBFhl2mWVXQdz25foHd12s8zCuX14MaIu
OWSk5pReyPUl09oR/eA9rHokrH7n93uTfB9Zky+OYIUGvpOeeZNSGMatSjai1uIh4RrY1RraBiGN
hgg+t70wAK57V2/6RxgIj9BkZWDUVnaSKd2MUkm5LuSCHAdSbq0+5MMAgAYIxArEuQTr0k82z4Bn
lk+T/tz3Eq1n+rfEONEx+NvtMgf4V6jIMl0RPYqzTsGNUMwtEYw8jGU14ub2KrmUe325jL6eIF9q
INCr7CX0VRlu/7qGfZ50RK87pni/HAC8IQ1V2eVuTL1eoY9CCXVL7FhWSCBRwD5NwY7GuEUKFVYX
8xJWc/Zy9rWzd+Zct7viAFW7k35Zo5VRqQa4NvFAzLXNV3Mx3z13Ql51fweg+HZ3FX3Nq/Kiyv1F
qLHnyUFw2sa8n3RFFHIME2Iapv8ZHNKqBwNnjGKcYBQdfJeS73EKhjcoWuUEbIk+F3IrnI6WUTDo
5iK9sf8JE3Gx1UIsvFBDz4CFWnQ3wAFaNctia4IQ8F5UBDNPrXid+dMbuMZ02V80JWdZRzycTm3T
7wajhNGCtqA5bVpEzcBmxsGRkhLZIAPPQ3ci4uxEEaqq9JS9GSdjwyHMJ1xrz+QomrJrooCjicSr
1Cx6aCfsjWvUuD8QjaGJFjuaOLTdEvr7pMUpjXZhiDWyynvyPW2fX7VJoyjWIlFDdwHb6JfGuwC1
K6k8CHi65kxvI+035rSZ70s/q4DIuYnhnadM+IFw21werG7lIBKDZdJERXNsGrMPK3gY3yc2s8DY
pGx6kqBKHdt4Z0RneCG07afrWiwIvb5nvdng9N1X+bQJRcGuKVExvVOurZXd8lkI/Kl6f18UW2Rv
Ok52NcVtAdLRYALSvgWzVCxUyaCjTOImdtMLSFIpyJetm2QnJL6DoeD6eQPTHgDndZ7W8xy+av1f
QbORqAkv0CZ08xhiYOI5YqAhnVGIUu9I1IDeU1xpK7advZTWornRJRo9jfYou45OfHGB3VusKkME
VZ8vsJx10RGCYuHb50paO9UkZbJwEN1soVeUwkNBnqoBvFL8KMDk/msSMRRYqnAdpR5LUW+PIU8h
gavAwq5A8oSWp9Mz7VrPhEXUSBHnJXplWurNmybYIkPgoGlZ2GNAnv/HifQNDSh4KfBTosPU8anr
n5b77wrYFVLf0CiKSbQZ0e1ENXlMXMl8WjHKLva8JzqGoXr5f+L0tJPnGQsafKa6L63wAUE6LWWv
1bAWcrcnLdMERMtkmJgMifGT6b5m8K7OMz+ytPXA7xTUMpJzJftiHvGj2sI5Kc5o1GcKg1gzTemp
qPgr+s1BZr7+ouba2YF85Bhoe3BEi8LGFdvcFIRP8CKVzp60EevuizBfbCMgQfrk0esCvObUiIKR
BBLjNweBe4hbr+a9kULB390jFFJ/BNTczjvZ3bX1qsKymR5lxJLMr4SAjPqLJ9cHQ90shWiNNDu9
NshSirM6Y/QmwBgR33kfnY5esCxCHtUOju0L+bOuv5dUz2RC6m0oGeirgFth9fG5/UOaKtquk9kN
l7QvQ/YWuSy1nkCrxMqgTKqXHWB6anTR6yL8SG+hecqyjsiESFME6bUAo8LY4fsOmwCDqicPWWCC
7ewg0331u+AKFTLNu8R0uRjtNbtuiH/HVYrdfDA1/hKbJpwecfnncxdCuEew3/XTgmssnvD8MD/C
tjlRhoXH/vQaNCsOZ3F0z2U+wZsRIiySLG4W2QZDx3tQedDGzr7ByiRvMrw4GLGyWrXJ9A0DTZ2k
JZEsRQCmVtfZugenquZ+b1NJrI+8N5oeMhbv3KBH4rDGOZZFBCp0p4vJZBu32r6U8msOP33irreK
99vztHijc7rCH5lOpdoJDaistKHtqV10dhEamO/hJixzsGr7/DbJpTEN1bPoIKYquN6JnlMyq04o
IPCCrhC7WzKFRnX6dYTZ58Hf0FEM2vqy6ugfenlL+Kjwt3VWsueeQedPl8YHF8xgeoC2UcOEG8Lt
o4Ah86DNAfL/ayX7qCM4FaVChtKVmdAb+s4kAszyfz7uu9MB/cm7jWa2RQWEhYHj3KGObaKiqmd0
1RbEAuMYxlEk2zdKrCFDuU62n7EoKfzMUUYHzyB2SL9bn9hDDNOgyE78eyezA26C1gTRip9IQ+CJ
1lq9i23dbXTEiEWwLyiMKY0ibJLRMmfglGoaL0JGdSM2YRpkpzz4quxbowekn9MhoR8zjkyPQGir
5MlNpArqGMChK+YoAKmh3TMuO7a9jxWY4fZHEJX645Ufvms9OSYb+GrIGDBb/n+JxnmyFEMhNs+O
A2P06DMtI5I0+TjmXY+o067tLgpGqmZeTvBOvsP9H2DRPhsUxysPkpBmjffdVH8WNUrSj618slhV
a6F+1eZIXJfHPHkN/SEcG/X4/33JdUn+xeVh2kR68ccvPX2okogssdSO0mfQ4ja7gB+didKkXJho
rw6Z1opeZgiiAv0nIX7Z2e0xGuxMvm2QSyfnBxSKI+Zp22m8qQNbAOZWqpKfToxKgK5dllsaMH8Y
ezKXZB4OODItN5nvgNYg2N2fJlmYhRYN0kfXHOXdq9D28LFHDrjhw7Kz1ACA7BjedD+e1e7uCg2j
6zTZR4kGZLpvPhqzKG5kHDICfQ9itnEHeZVzJNchHLCaMGT9Y8u9G7VpSnaTHz7NO2IU/H/JJ1cz
DFYF6n5Eo2S9x6gRhBzjFvg7AURByxcYENqs8b1HayZZ8qVhKZ9fWydF9KD+SpvAFCyTw7fCW6M1
HvW1KLssIFE7Qme+gFuxdD/cmqZIa/HMBm0R+UU5lsUfINwkpXNG6bVkdcRLVDj5nitZQavZv4kO
nxfqjW8UuSSh9TkRn7o2gln/nqD3p0g5Mwmr87eDypk7qGmgM0m7GoezFVPqxXdeRT4Xa7M1Lbyz
u2+IGTvCHjv/MW5ePsAH4xez8NfjlxwpmY0/kp5ZYrZJF6pYIyAz3DhMYh07dwrUeejSXtbFcBvV
vO9fd1tWa15BfOc6cILDTkBfBIehNstzDjPacIfwBEUhC1XB08sJzt1dhx0MW02/eNwpyH8GGmE8
eLIxXzuOdJKn/Lb+WXSXvnW1+T4ENqYllS+Pgle2Km264+OQl3tmiYYgmrj9lz8vRexEGcwIdLrb
akTEQLiyklMX8rVSLppoaKWGCgWPiTgpQQlIOrUrkDx9y1yJmewVYdEcb9UWxhEdXFJ0xFXD4gUh
WkhMzUViEGeaTzqL4ONU6h6HyvADWOH8n0N12EPFZBHJId7TTWDSh+AAM5lxbwKnqN9X2mNiodBE
4hQw9lDqUR7wuJaHArwN3PqcjJ9ksyymnfd8desbh8KKWcBPxbv3rRN3iQzv7Lo9UBXonqt17NbD
TgVqdmD2lVqR8bODOVLZqUPoqBIObe80F6VEONsXGTiJMeVrg8eB+iiWTTzz5V0yU1UinSUYkePY
yAayTdwPRUyDSA4Dekrns3G2C4L53Kho9AjihxXtVD+i5J2RVy10ZXGNgUbG1Pq0LGsXyYaVUFcD
V4YTSvXNUS0saQaBI4C1Frn+p/kv+rj04McYs3lVPAs17jnm0KsDeFOKTxscgbF+axqyYEHXOEUO
aGuyVMDiFCNuzsifIlDouvcB4xu9LSksb3va1QUJFrU/unv//OLL6H67TK0e0MVbiKe6cj3gKgBd
ZrNGEcM0myu0saj6pl+lg/mwkOTi1OHbE2LdBxJauCeU3KPqfvx7wPbttTYax0IGqaitLn78Lj19
fw5CDDktTShNRP36UeaF/UXXEDbmZmziqc06BF1wudXXG/BxOVQRvP5F4EQ0/sw2fkPSMTElw3/f
AxPmUml1480ZWdLZvuvUYGAHoQ+vaNJmFaf9U1mkgGHynE5Jf49D+24JAfSos3DdU2MpNK0/qc9k
mFsxp/qikuNU0bSkkCx61KL0qw5ZizT9uxc858l2+AOTkz3pSnEQT6xcAiRjOztFSsyPPZRB7zPB
9jDfJnRI7Gga1/Q6OhrE1DsdRa6rVpoHfPeuAfw/d4WnP9YdFDnkyOOI//LCnADyp2P9J433Vwb4
SsktdSZuEtPp4U/WUeA6WbWIqI7+A1FVOgYF1tPqH4R8y4vYXE3VbNNh3h3nrbTle6QpUGh8qFh7
v9D1aY0C7gLCGImzOrhB6lBeH8H2q1FJiowpijnv7uZIccR1M1ZsA5UChwmTvAGG72F+69GIvFC9
60oLcQ3xEF3ELuJHYX05A0qVY2kQTr/Vg7oKNfxPf+GLE0z2uhMucda5uMcy6gcGE1nBSvK7DMu2
2UJi3b7hnEBsotfynQwgHfs2/Lc+TbgiV8TYi8TJJdGB/vPSjj6COalXCzFHp3WY8vv+h6/i8KYf
bp/Vv/MUghWnI57hHpWH+DNLkIgAIHPlRiEjIGenEchMP2j2107D8n7RPcrpCx75urO1djz559Zb
8cWqW0zRI1Eu04740SLsmc7hixzyqomIauIuiXzd3KZttLjUfcen5T4Bx9jQ+ZMDzjgTdyi3TS2V
0ib12geUhNxp+RfFQVOvCGU7UcIGWULFlNfnsX7cQ+C3MEsJbPGsmpuJVDWUG4rKTv7mXcdgUutp
ybJWgFl9FoWiWZJkpaQsNKSULohNqsRkp+4tnwiN3zGUXBN2ogNE8zkwD8JhEFjoiOGmoCTDeDYK
gKN2xDL8To763QxmDBFxAGNro/jIPaHdLY+wzlqA/vwXBZwJUHl8f8+PPgl/iNOfRtEevKM8Duf8
h12/Yb+pvbU8mv+kyUSOhWe0hILRwu51qE+EA24MlphxMbJvQLJh5iuEoJoheBeB61hzo+2tJJiP
IY0PCu1q76miiIdFiNm7ghr9aQcdYTHgyx0r1+pZKU7UmvJBZWw+ElnHLQnSow4sG7TJPLmt6USX
fiqHbIX2LF5zBfjowDREKkyOc+xxUTeXd0zDLlr7JZauKybt2IPEvl40CbtslE4i1M+8vVdXN4VQ
ZY7+ATsUoeBtiZvTDuLzwFIFeUIkfpbzhzEpppdS4kByVhHrrV1kCSfvz48CQbiPJaicluWhwZAK
NCm7e6UKtYyPTBEB+HFNTxEfqX+dB9/6E7+by4OuDYrNrAGIU2EXBgb+Bf7mGkkXr7+fVFdktH9X
u4Hb9VwIrihyeyPs4pXKgRoEWwXGfF8MHgZ/GcIG1iEcoedr+Z7E1f1TZtB+rCZExs7S1uaaXQR2
Xlb8TP+iokv9x2NBAeDvnTwwtpA+bDc77Y5zXdRYPp3D49N2fJk8bH1K4SAUdMMrY27FaS+PrOiw
76GSuWr59YViPV9I5Vz7e2v/Mc+hcMVZEE+teSjC/5b6YKo/0w4QDTqbZYgcE97FqixUVKS2q5kF
PhZOdGk9asidEhI++O8Rgl2rQpatLC72DmvPnuJ8Wl+qqu0C7qviIsjhkFjdONb4xGr3kr+wbjln
LQ5NMOOIvGUeVp7UdVF8jrFunAQ/a6CZnhPdx9Vjt/lhEgAxVrLcHxOfCDAATQXasSrB3Bsu8Mys
x262txiMlTG+GpkvQmq6vH+6aX5mIQIRuZYYmvxewjB+LaP43l6OXsNsfiuhCNNj1xwJ/yrAUyna
tQBhgM53WZ5pEGsPjudQWiGX5sGRmyqHX9v84fN9i1n8SJqvP4SMCaKqNr68pISvfXzLcxHq8BW1
Di+UT0UKoibJ7E8y2hz38Qu9Rr/Jvf2fs7qRY/V9WL5XOMIGE3Q/+pGsS5fc8JeFt35rVW6WZ4zg
dz3rkSiZS4pDk/oHhBkqfjqFSO4QGhYgDhjBpqPFAKZhbJwo4ZeUxG1Coa3trACZjtc746LDLh1J
HEYHEOBSec10Hnuyec0xeul1vKm4oBGyLul6icU9sVqvbbk8/mdi4yDo+9Fx+cavUf1VZ1fh1XnD
uPUoBfK/vE/yvOj5G4wazGIjT5/K/QZQjwssgk9fy+KaDlQXZ4iPlVo8M+3f3cDc7HxkYYqy/7DZ
033LC6FLFaK3Rfg57Cexv06Fm8vCbyfNFqlZYmHzXloa2fFY1Jg5/rzP9QiDiYSoNVHv4toXross
jPK5DWdse/nTonuArI4c3olKXeVNKbHtRrt+eiqMbpQMSK03BjZdKjd2WcTsVKkVSsV0azQWuKmq
t2J6JXpX1cKvgyNsNni7hqyUJELN/2Jcl/ON+1u52ErEW/hLEJtONxFu4/M/H9c5hh0BEIDxufaX
k545im1I0Pmo4e/TSqEiZZheVNLY3UCi3ukQ+Fsnu/3KrmpTywN+qTHuM1jz2CPm3Jow5ksj2Z3X
5nLsvF2PfO4LEfjNWJSYp7zMl/+o0iVJLv/4jNJmxwXbOZ7Qk8vzPWBbB9yyRMcJGv7N/QJ+TLfO
W2KeqcjukaoFqwRPjEqJgmXm32vvDFCqeauSqU8mE4naCt3AXtxzSWstTrHvogCGUA4iVigkkCDF
L2XnCnxbEPWdKbd+OXg6uFEiRCEaCLzKwaTOoHMJk/ps63kqUHIaJDP9YalDTNWg1RRU0TpBf9dN
XQbwHB8WEjTDHJEANR4BHdX49j4ZSVhIGup99+CglAsqRHrZbrjweuY187bEAdGWMoTUHEHEVtuj
m6aGhRi8e81rPdWayx/xyutJf416dITx2lGBhd0mufIx19lsdNIN57roJ8K3hzVWSoTzZXir+ODw
QpBOt4feppKLZRPA4SFlsR2oghYW2SOIs4UH3pGA1pNI5I0SNj5+NVVMf8+AnOnRNd3elTpfmmT8
2+RpwkjPYtt7/Gg40enm25CFzK47kBI8PmagD4Apox4NV7GXoY7ClS2gn2ibtzTHPBpBaJTPU6ma
Yc+cXkydtxU728rKLX+z//9eqwONCS07dxKfEnOUpwgtwtEO65puRRrn6nNcnILH4PMHgqOY0u9+
/u1WyW+53OUw9Wi6vQGZY1RQH0tHU7MEukoB01MssD4HNfsSu2iGuwfQl6pFZpqHa7FQklyQQaCi
YcKRqy5jWLbl7cFveOfKNesowrJYA9qLuo1tCP/IgoFca20y0k3GJdLwbF/9YVvJAGnrS5VxFxSA
Y6OzQVCPR1aE9ty+w7iQ0uNcFTgEfVjhdKAcNByNQcmH4gahEPqbkCLkPN1tMCp1+MIOrLYrC7Vl
6iw9TQGsDfzB1Njxz56pg3uwrePoCI24SY+JI2ZKpaOFJi4TkE3vv6PT8p/ya1jBvgzVecVL3Oml
PC5TRhVqEatGISIGu1Q5chHDNg0YpRjo16TGU8YKavVMkVCpK5+wvo3zRkEEriQhAhJfrpP6y660
Qc3WxyJ9yzRZRjLq1jMXr1MmNQ1tZnFYPDpVPFuu/hOMhFw/PuNmLdm8CCv5B+kTUeSf8jGNu/5f
gPWSxqPbwFdhrWRW7k6i5EPDExRBK9oB3IorJ6idL5YtmZAwMyvmShWRc+WzF/MEDoupIQS9TdWM
o1FB7LCNM8N++iyVrbxuEnN7PC15oAMj7QbtyJ2B+qbE489Xy3OIo/e289HkoQSUhTOdbQ5B1kwZ
fmjG4cMau+aheL0BJ67kcyHv9FHPon0H58MvuiIDYKwoLLH+YSEMRaHdEh5p+hGt8ycNt/guJ/dg
+Rna99JPOZS6RymW3iL6ZjNiEvcadJJshTr3V/O0YKCH9DeBHlcl5JefdVvr0aMcN4aU8juUAfZ4
dGYtbYM3RipZyHupHZDOLfeM1zmQRisOS16K84KRHrXk5kmarYsFunbmyaaJoJPIxs/BqMMsy2VX
NbBN0fNbxc3C1T7fMFQtS139Y60CbERHCJFxID9WsNPAnTr9ChXkl6u8zkdI1QVWS6cTDhVSFwgV
WpMl1x/cPwIfNtKt1vAsU+Ft/P6IKfJvMRgG1ZKzb3lDaGuD4uHCVE+GBpEy1RTVipTRhGBnh3BJ
wFBzs+BJ3Vj/EOZx8uKcz/fymR8bW7kmxqc9F/Wl6KtKhWgRzKZnJVLaCSJ9Zq7KJPvM4wS6K1fI
s7EBGexw69whCZZ0fqoAVpSS0XYgRkf330fggllC3LqvwEt3bBuII9SouX7DBzgKfZs4KkJAcsXo
A1YBEMCDVzWGp8chbz5iKuBFE0I/rG++D7wEGgHtF5Sl71IWCDVReT2nw5skf8FBWYDhAzjTv6wT
qdbyVf6W6wt0m2kJ+DqnlaNclBVXQZZ5WUdvfSslo04IJOW+9fUq5k04xjdaaKfJN2Xi3JK6nI93
bx323dmXcJQs/xYC6rQPtoFgGlu8Ufqxk4XICNr5INGNTKFFH2zHdneQcCN3wnSpBeqWYkYZZrKW
+orFthjuqVxIJPc4GTDdg5n7cV4jRotgu+V9Ad8fAoZaZDteMRaUK6hGMVgwlTdLPj7gJoc212um
GMuGYV7Iwap/mDDOQkye/4w3N74q+etQv8DbT6L8aWdgfQm9mxueVqkGtNypNOXO+E4oyTgc0lNR
/KUW8DAPc+yd7vNK4kQcx9RKeBb9Bc6eE70qbTMdHwqldKI9ol73hAnhZRUi6IBGxjbxcWgoBT7n
oZ8Gd/4w4upqFLgzmDsWrhzWhVf/XIAGe4QpjiWeIG23pvSWhwYY0H7YnTPlVNCmA9M2EMHPqgGE
d88ndaoMJTqmlnxMkQB6Lctz5fxm6H10d2bfQltqH737Ngx8MRXysQD4Pf/bgMr2pmQPvCEnbHpa
bRWnVc17H1raW2tk1IP4ybH1hE1AopBAr8sEV7MfuI2Dh2RpVhPYXoUnv6ZAtGPu2AcdC0VU+t+d
5fLmtEHjnPyambcwLqeGOqLkWa2bsDEqdezIUC6MMazBeR40NrODiadYZx6MoPXp6SXI+eHP0Kxi
BaMaqa0r8uUGcSeSTr6XU8n0xYwef3tjnTdHKvXVOdE/6aVmPOp2TDKvdinK6E9C602mMXMv2Wpp
R3RKtNS82YOWm4+ztqtV87sfKCP2Py1te8BMhOyiVKbALD8/49AlZz4Riu6e4vTmp4X27ILJpnEm
+oe8ZGR/bPeDyO3NBFGwAywm4A4OLuwx/KZtfF5AdD6QTxE42yJtlyGpb/aH54yp23Op5bVHwWrZ
W7tQ7O5qRFBOi1H7rFOJSx8Xwk0Em7lG505NIJ/gM0UvIhW3lllR7WXhI05tS+jCNAw3dNQ130CA
ngD+lK1ecpuFvGLf7/mzERWSIMxxCEdmrPz3GtwddXl9CX2NyUclZD3M3FN8O+31aqmv2xEWiYn2
eSDVSqHQgq9YpnA0P6Iw3CglImcLnpkwO6SZxkwZIfMHNZovNwsN/UmgOEUJDioYb6dju5+IBr3S
M8WCcCi3r+RwBUlB3VFJhrxH19yDMxqh/oQC+rHBSSPQUaaUTzzbzK20f3viW6PCoSszSMFUMHym
ECI/XkpuBSh3jCgqykamW6CsTYXRDdSglmxgEz/ysvNvGLPqisuGuWO+EFYPmWFL0erKZw87JigI
vnrY6zXowFhwWYd7GKl/GDgB1TPGMIx2qvWeajGQfv4jip+wPvlVzZBcG3zgq/YBk97QdFvhxMAc
bIE9vX1maHgqpSS0gxDuLCHLa7GMB7LRYP9eAEal2I+n4kdt4gT9/HHwESEjrJVx0W/sWwF8m5CB
tQaOErr4QjOoiVlEIXFdOczj6tWEGlDcJwcnpsqsiX6vXZHRAR/xFOSxSLokEo7qBr+D/NHOphUK
VYuKvm+yNG5iXNpn1TftdV2Aj3k1UO8AVeAN1oAkjji9hSsdASVCgVbljuJYc0pwSG6ibXI641fl
njp8OsYzt+1Sw8Nq8qf5ErXYdECad8tlHOVaZDW4iZSbZHFChcZHvGzPZbqGuZZ7rT3mdl/h6Pdx
UBICTXiaRfmIkxs++sVwBTzYq5iR7CDl+0NwP01iDXxV+YrRuDYolMRAA3ZjYpquWrxEyuu7TKTV
0M/KhjiKTYzXJy7nG4TawcgA7Y+/ZBk0P7StDgP7Uwsk4D6gMnY8MAc53j332Q19ySNBnzeZbjAi
x9MivgJU/sT6sy5nzUx/VtUUoPYNaQAVj6oqpW0ZR8kE/NHGNaXDnvI7yibNE9XeOSOiHe283DAu
rCFkUjRhlJ3bKuu1L5YVoLzY/B/Gm6CDgj9fdCa0UPX2+crAeZf/POa4kvqVWGEMSfM035B4zbat
B+2ds5UDpxqyE7kfu7DXp918VVWTqph7leN73xQY8d1QCRQjWoWApDbWnBRf+VuUJ0Ijx3DK8aWG
W/vld20Rvvz9ZISPwQ9O3Vz6sOvTwIbFpAaMTgZBQU8dS1JHYj8P8UE4l02a++HwF2Ydxje5JKRG
H/Voi2PxEWrzrKx73u6n38HQJb+wyQN+yVvd7zrX4AKTFpaX3NS/YP/sK1p2haPOA0sClABBWGJH
ky9q5tl8BEMxKhg2NhMpjVW8IU3R93NCYtHoyXXLetlyJynhyV6elU33x2RKCC51kZFtmdwpLsNv
u1xsRao+aJAg7gQVCb5DUR0HFjaHJCn/bVXhsRL8z2jrRTJMVEhLLEQyIvxEHIMiJvmSt5Q+BLNG
DcWfJRmxm4FCDbwmjRszjGKX2bVm/rFyU1S4Ef2uLa24DxivwXMtxzUVZcMF0RwJ7fn9ucRlfvAL
1gRIcuAI2nZIYKR1vaRfUE1i55JS9AF5f5+grIjPkLsE8Uvi7gFYmWqHv7iycuUkQff/mmmpTp7q
sECu8AehRlBZt5VEQZIXd+4s/WXExnYEt4hloAaUfwkoM0LoJ7YkhzDeqe4S2zAn/zfU/r+mniAg
R32iq4tCvvDH65bdlvN8FsterKncR1nqDlVbgkzRgGZbXlBb85THzbPRsFDSvP17urjKmC+ePKvu
GlYGrrmG0wxjI2x3bA4Re3HvJN8+yLSBM8SJZmx7KdRX0DC1xsEo/aWkRC5t4XfXhY38QUtPD7ty
VlHjaEGx99USAOCrELku5T4K/j7GZpk4sWGspcbQcA7cSNIrEyjiznbvngYbErXmYqj/Ub153jN3
wyGnWvDxQCqfUwsSllskfyFMM/Zxu+/dN9CMvjKbH+ecRBkgezodIvxZQ0M0hkDTEQLeOTzGtSWC
gWOgWFsOxl34bUClA6B7pHXMgntMZp1nVWhoEH+T0ib9nAPG2iWiCW96O3CIvak02znzw2odb2er
6tDxFgRA6rlZ5t0Rf3zH4V8f5PZroOjoynCDWyuY2eDIxlxXfucRFNXUhxMloRqQ/allTXqIfawo
9/Qcr+abdtPIyk2AYx2BEM3NedNP+jRZHBWWvrRCztp9Drrno9+jo6JT1Gy/IwpSPszz1pA2JBzF
ETmAgb2mWdMrj8muFKL3Dbw+ywGzxFmBUhfI0bZ8j0MCiKqXDqHYoaOib61HXvNMuQ7Kt4rAy1f6
bO7HMsnCDIICNtucJrzGYf4Tg9Swgw3DGAsdhD7l7y4/ODWKJN5SGeMiPbr+TGVX6Z0f1K9qH8Je
ARluYikhzSZYTLNA49n9uARmtpjMtPrawcajaOS74HbNSH3R3k59qSIkQN3aayeB8PXZ92htm/Ag
gFYtutLoG4d34uNNwhdZRBOMexG5ei6uv1+3yuzK9JrnQkTIB/APAz4PDxKnzSmSfg0VeEdix4BG
RzYZes5AiRIHKhxepjfZAZNRzwvbq/7jk7Kdz5XSIHLGwtVaQ1bzu8D+tOVwDNyjYX5szyCVcQRx
lssTYQZWro1A5830dbAKkmAfnxrJUW7Yd5haLYvl1RCgEe8e+Moridofw2CDNT4mp89e77Cxb3yy
at+FAhPg2FqkDWo1IlS0ODdObD8KbgG5J6mTaCnDJ2uLWQ3NAznZS0lz1Q6vg1bxCRW9jEKjuGfM
vj/u8aYmEEgNx7us15pArsqr3USnCtrhFo3pCLLstw43bXPDU60Ged27kmb+tsic9n2y+wg/raDs
JAC7RmVoJD6GoVHmX+G3lMu/45zZvL1k9O1GM90g0sp8/E+GFftdQdJ1zf50EyL5rawVM67VhuT+
yj3hCveSvIMFRVbXpiYDpwyCHT7GGKX6EMFUt8ZEKlCZF0GkNG4nHzLrHHtBMMaNqKWbGN1+NYXX
nMbfr6+1Ah2bFZYHIXRYYQCznXSa5Lb8XjIWAJlJeE1syio6S+XCnxe8weQ05mpO/Gi+H7Tediel
bnA5PXIkS01v7h1Fh/TlSd89wo6ayJp8wPMkPw4CKMFkgCfEpBpMOUPSap6LLVSvG03e3idw5qlZ
G0MNiXzjfaGWjm/+pZ/W+0UycA59LsAIWHJugSPnkvN+Mn4zA2WJqfodsuD8JAloTn9/pA76On7a
GcwjML2Qu9B0C0ZFm3+8kSvVDjG/SYkK/2x4XWeLfgXsMkhbAAXM2yBu9pS7vWwW3Y22tfpxO6gr
kVxV/UpDaVkz+EtMkcJYSU6fvtDFqC/y5mcE+pRycEmTGREltX2WaDHt3AAf83R6hZo6eyLsum4H
k7aUKYNDVnkHbJgN0SoXmwbu5il0ON3ec7HtAghDwtnXKBoZmO9868Ks2RM/4WQpnXyk62oksY++
CBcKzrCySWuDmLZnbEHYPjOaJGlKSZOUU8LhTftOM8Ev/3MkTF2qfrG3y4OqEIctvz79x3rM9u5n
4wtrjFqCRZoHHyv8mICACGkZ7+UDxMnntJ0UlaOah8T4exScJ3soZXkfJaOCxT2Aosm/O93iDkDi
Mr40Z/J/x6x5q/dvxPJkTZxBwvyYhvjlhi51rY1pjltx5oKxnERH9NPvoZf2MSfJqQQFBlbSwVFh
FVRyLYAsrJUsruRiI6yde7X+uz/elbEfqif04KGE0nAq5iMS7g+3JSy2mworNgV6CLTgI2WSkxng
HqWmakpQJIodAgpovIhgoFrs9vakjNaH/6ak2kQVU1HsZGqJJpTNvJmRUzeZSldRCj1E2fGcM0N2
yDeu5SXMBTMhG2i8ECMwJ3LJP/JUzPcdVjtF8QbXaST8sS5cq1dsYhgfRoGZpivTlSDNKDiuEEVk
QGpaNBx69vJdYD/ry1bGrgFWTP3HgHbHp20lpkwvoWH/oCsjG0j10rzqLyYALTxN40zOPsZylHid
NyyPnOt5skAVaoEoei7kVc+Nu5O18jvZuPYAg/uKA36DGc0Qismnoo35Gbvmxq4S4QUzvIg8GGXB
9I371v0j7iyGXkRTQclTNTAhSHOFXDTXnAVLcQPUPyFNFEWwFJcEN8gvithj2HXD24nYj3d6SCNY
d/kI9DhxA4Swslj8oMXauWkq3iqJW4bS+w1w3aIoI8hIu2yGaULlSNFrXe1HTDYRGoVtsgOCb+HK
G+gZN2+EYcjX8wLEfZ+D9UNmMZnX6U2JL/AS09VnYwsxR5UmJ69i/pH8sWHjhCYSb00a2FWamRe0
F4/9qbaXJLHYfSKVa/aQ7QxT2mKLgyWz8OLURhXMXQAkGOhdi2JWLboahx0M5HL+pu/aMyScDPk/
3iSWZWbS7KGPwORQOxAIqMmTwqtw+JtIp8U2KfpnGHsefLJQd4UQj/CVE1SpU+htcDRVs4yTpb7T
Ephgdh6+yazQ5pcTxQADm2PJam2b+LrugEJVjOV7TBPnD0SPNTDMG9SUdDG5EcdNzGGv+49VTtME
kY9gcbTCYT0DCj7tlWCvTlev6j07WF3wEvj0d62cP/obEy5lUhTmYENvAoimFGZsAubEJfuG1M4j
zQyleLGUQFoc1vBbQY56RwQEomIi2h/adsamKuFv5WB3H8OWmwSnn4w28gy6APxNARINC8SNqZYq
R1NkHORCweg1Bn2tcih3RDz6RUfKQP0oV+7UF2HFmOa2/ZlroMMrK+NyXpLbdR7bxNd9WgWNBKz7
salXlkXVhl5P7FktDFDf00CYBk2dUbyWByirt6SaWSLH89f/ucJSrzLBK2VJU7KcLozbhXDpzctb
4yMsIBC318RMVQSuy5HQJz+BKSHow43S3Hlj36N7isyrL+4gA31KfwKX8TByoXFxvm2gTc6EDv7M
Dwv6YlIBElRDcClTx9NKWAwKM65zMhpOclLtsyyLAIP6OTRtTXK47Te+kL9tE1kP/y6I7AN3mszJ
Pei7gdIafhNhjfONTQzXO1MD/emgFTZ8KN1gRQF1g3ep37YRgX0+nexdKJhQtS4m1QGIQPJmMb6V
mSepej65FQV3iVIq9rb0L4OBU9rzr9Bes3oplawH/TDV8ddiqmmNBYU5slnn1cY/C9+TUwPBruRW
sxrwlnA3pshkAt+EypOvmQayacYMmOyRU6EeL/tT9F4sQZckj6mzCAb49uRXSg+iIQuTdNEQyREX
lm9EDuDbbzadCGw2wN8XrbffeVNjzO8zU+PlS6KSCK50iLhewK+4ydvBa3RfEmpvjHVoXDU7VN1b
AmD28kOs/ypkLroxaw81Dwrm/PLgly2N+NAvsHPhZwJactqwK3IlZW0PzBx8r61XwXAjSlWabwQd
kqAcAirX/W8jsV1Izb2jr/RTmho/2OsEiVGujChGjwLmXmnryT5nr22WF0TbOXZRN5/ZC6mQRJqT
rgRiUytmF0cK6kuBJm9FYYhAyS6RpFUx78lN9e0NBnW1ynC3QVNKamFJuK9ZN7c1KyxLs0rA4zqv
Sekc/BxxF4AVjVmu/8pqcZzdwr1XqrBWMuM04stEnM+JWu5TElnR4o8TTf17iiNK/HUli4x7B5Cc
J93SzIDHtDIGzGGSC2Lr2aRGxkKURuj47f+GGPB06KMV4Bu2ZMA15HsoZByZurIBsm9NwPYJ2hiT
ZpCgAErB/jA5Lol/b/fcqyoHc0GVIotyYQT1WB2MIZep4iMLSclrb4hRwyq9v+4V2eFonm/20P1N
JqbbSg8msSHmp4sSs28fquO7/izCKrapbg9tfQGeUH4SwlvdLdG56TkQ1ZseFnbVIJyuA4H/DWQr
zsquIF/9soGjy3kmrv9utpzGAMEGSmU0uWar80SuUcS8rqFeo6FTyRpDwdFqetIlVS9UBCobVTN/
G9y2dNuEoGFvJvBLSG/G7c6Mxp8/yqYte8Jf/Wx8Ad6ZXF4qZugQS6mN/riAGvhQ4vtB44yadWcD
ivMBleBgKolAvlynJFRCN5Giqw5SgjTM//UjJNxx7X6Xc4U5tF0NBEGcwxrpm/vrADmVt7oCHX9j
gZD/6DhgbsfHP+qNyrHdSLqVbbyu9YMpOP9poZKzJX2EygdmXRhQWev5ENTHNgXWT2nR2ikhBbt8
fHQhIScbq+Y43Q8852X4SSXD8LMEWMBfvWtZUkMPY2JPnDZaR59nuhtu4fBJZodMrf5cHVCU5j9N
Pj9LgUZNChmM076ybFdlWrplqPQ2LK7fZ5e91EA24+g5d2cPIizKgl2Cgt+Dv8oHPHYEPhUCQ8jM
zez/AUZcLhnrYyuvfBG0npCgpXQmw2DTr2QoMI6/PgPdCxbYO/vYA/75AdyZPuR+Vyhp7IvWO8DZ
XS/terFLLuk3BWmXCmbNAohrOI+aW+Wf1crVmhoICZn6GB3vQDn9rJv0wXUbn916PWJf3vQrgPcQ
OF59+9tZDQNt3VcGOBjz05l+w50L1Sv25muMhNFmJWl1X+xdnOyG2yGaLMCtkEnvvERD7+lyhAX8
Kve1Logw12IvUxjxEy23fTYUHCKFfX4b7h6jrlS3XXhv/txHg8G4d7niss8KaSwJe0/2IOteEET2
nqBNk+HIssUKnmYj9YMcN9kA6lOvwqrKirDgMOWDGv5KvQgNKF5O6h3XR4Viz6ZYIZzIMnO8XKOQ
Iv1I0D48W1UwmSgpFwrgT1TTxicmIv/TUigUWjSnz7UlxbFkAr3BaIh4Qm9vJwGwczDqfnAoWowB
oVMjxoCq1LuMgsi9hOsCWnXuq/Osmuo3OwW4p1ScJRIOlcHb/oXj6pp3SnZb8Da7SxNFLIaX/NkM
p06yeACHIpaBYLg78iQrmiSIeJ42KL2q59aJV/pjomqlChx4RoZ+qC3lgjEx0FFHH7CcxE87qfhc
Vo2OAxw0TvRuJG5hQYRF8JQsU6PRV9Fh57rAAxVP/ehWU7E6HHgcOogrwyM2XDORprR/Jo8i4rE5
xQdlaC27oPpv6Dvn6dF4wwluIFglQiZ9kX8XoqtuNvrjLBWBvt7SLyeAKtS6rnN0JmSaNuqQNwVx
YLXFyXOZPyXNITqS1ScH4wrkf3irLgvTyX2+aC9TDNfFd83tJrno8ybFuXDYediBtFGoToyAHw50
5nFIA8+GG3pGbmewapZ/ogodGc/2iCDOD9Fi8hWsm9tb/0Ouo+INo3uVRjrCxB5rHTccFryL1tk8
ZTr2qopgW1WOrGPyLQs7bfGfm+fBWQHhuCvuqT25dh4SqCFUud56uLErENww70GCqe+0tlzIjKbH
6tziMZb6HV5aKRPRNYe3f3h7fuzNG0h/cOqyZSZ8qRd8qU87TKOJSn0FFzI8NFv2qDUiUDR0tvCm
M3SY7PpIU72Jf91Gp1DN97iWabcsyxg26hPQkXXEWZWBY4P66BYyzLJJOvk7b/J8ODQ2Quiq/6MZ
imKGJqAZQNTaJgtLDPgtjCIZzd4fU/p4aULLpR1jMBBYSxSrBMXvm3mnL7rt1wVoi9CviI0Y/Xxt
qIybmOwzKERmzbN1MlvCO1HE7/o91C/iCXgOFjYNq/kDuqad8QnAg+oQE96AUQqW7frgxwSh3LLA
C+GJPFPc6QebPxGrX/Sy9hz5P7mT+Kp0kf/x7TQiomXHqXCsIrmMN6MRZt0ew3Y5Bwctfd5HMskU
P4qj1zl8+at0qsiw5620B0FRPD+uBze+ZkISO51Savxlt8eOeF6oiwzZzOQ/zmBZrn4EYBMMbqCv
wpLt8QIg8oLXspOQwjgqRrNS79rDFH0b6c4i0W2xSm36dR+UiQWVJf3tmR7S9bcibWj1ANHg0ePU
WXGnKW31o7Qerm8exD7t4dk+tN+j4sDZ9tR0/n7NRZRzduJB4e77nlFA+phQfXBaR1xTCELTyRpO
IAqKa8sEY4XxFNV4ZTbLB/euaYV9ptzmlJBFbOUSxBYqL0ud53WmA+2T5KyhtTGdMaFM2x2IlsVU
J2DiTh8JxTwkv1BuPIQGuDnD3ntPoQvgW87fdoDyHyoychmveHK/PpLxO9kjVfs2z29fnfCMpXjg
a3qdsYNJrD5uODBl+ZA5PLoIYFpoXNLWLabgfb/dTJ0fS+eYrZcBgSCLI7pJt9ICZnWarmHHlLM6
+/AkTCFbtQX3AH3dAw6gUTH4AYoC+ZV2Qm7r8fa16cE8v78+7hEdiApNzJs7ehRUyLAlKy0VvZtt
NVHEWxR9sCyKJONbrxFyc5vX+abitp9jNRmdaUopDSPy8GxygbAKwPs7GCb4EWVOHpB9QwMEXgIp
D29aMH8dQnLotwaivRSEFp4qWV5S4mYp0lGSJnN01fLsdXZZeTS1Wp5LKj3Pov1a4s4MaMKLMNEe
hgu5Y/i5yRgItcEIE6gsRy6YYYfMOln23eunMFLjDTyrlC541pBDAhlsxNT6WgmCtJpzRN+wEuNq
gf1PJ1cFcPQGBLoQUgMY+2N34C8awPV/EU0fkk/BeG8M2ALvN9SOEYw8LCsRdlh3xTm26ZBrl+oe
gkCzgWovZ2PdT/tEEXkJb4ovNc0caIxm+nFoY5myK8Mmrn253ntuuMI9wyt9gE5Hg0ZdQ0OEPBz1
UsdbGK4lp0JmnZ5WT5nnj0FLRNxHelwIPD6pGA1eE8eycZ/elgDmmNPhI4gglCyC+IO/DmTRzZ0i
H74D7SpEJcMQdne8TOMv/COl79CqeFQ+NCXiCHwJD77Fj/mVA2/Qd5WFYcOoLG4iYiIfbRwY03C+
ek6FWSwVZD4KHezXdHs8hz+SkYzjvNN4ituYG08tBlvaTd4PYTWgkRE4mAcktsJlUfBRD4HkgHSt
BoAE7pAaDHYgL6xrCXcUqrJgvB80alKs3L1K7xMYWNaNKvbubZ2cKMNXDr6hLDgZdjX1Ng3a2mvI
luHjMIfBMGV5Ylae/pHKBSIXTP27vVKNdDxRfJkPWvLlzWYhI2MtpuBMe3yFGujeNYB+b6LrPJjR
fkH7oJhomwlBDaq7xto7S9fp8zUzaiOM1fBY/EL74PuT5EJUGkiC1/uzAHWpTPzNHlCKsT8UeVXD
U/wvSb1hCdESgxU2oBqPlC+SHqo0bFzq8/2n9TnW8+6+3DeGE8qT3yVm7CjwxNtjqGa26JWAFIa/
AcjT9BzDmR4i8wj80wUHWsQDa0lJg9X9yVuVMMTxxufLUI7W3eNLaiyj19eZANnCx34lT9pwZ0uJ
XbE0hv+ISgJUTwoo93nEceYWje+TtoXUVj98TU2uuSuHzHYijWsZ7fepLogXq065Ex6xmLV/785W
yQtWGO5qjEu6s2lpFNTv7uR4gI2s2WVOcGqli5aV2lR/rdZOKu+1JFp89ZCwtHZZ438J2BKSFFzk
tXqbhmyZ7H6oUmcPtuobhIzhb0mTnnj2r1X/98T/T/YnK4vWA7iHLk6ykkBV4YQpNQFXgQkluhRV
s/Z6iqWXubxNSAxuF9833x0oHjnxxYqN7sl0x88LedDSWhfPxtolWjpLzKiM+KJsMGdrz9/xBg5V
u3cxZtexIdf0wcRTgCioByJ5XeRWZ+Lp20h1it11lwHWvj1/7NyRdtZt4qztZ1pJuDsLKgufz46I
qEdjCNFtXymC5vmVIqlsY9pzorJluHG/eNJKsD26n0uCrSHjiod31g2nWpR9uUbCp/4DLN3F6srF
WQ5jregq7q4cJQZfscp2sToRt1FtLvEqSPVsNP/YGxs8tpOzVFSWTZGlMbttpATN5EP8O2IAMU0f
upbnNEI6lZzF/Lj1snmKc3vIXxTLYwU8qHajnarmWDbYDdhW63CnXyZGb8HX7KpVpChlvlXv0oKW
NjC721FTYV3VREKzwrP7/qU+Z7dXBUYMy7iod524vvFCl/pQCHxnSjjrUNzwTm6CfgiBYNXMelBz
fANwsLlEEqD3bApSD8jlszIaQXFSZoDOeRgl/cSe/PfyV6RvUO6OqaE4Md354scYTOCtaknzYEUj
HPOLRnVBGMUc1VT9redx+y02zphoULLPHetmBiKyw4xSnRNrU+++s8gfey/DN9VukFBxLiv7l82F
hJ7C4pv7mfrJsnRDWLXr3D47w5HYlZw0qm4r0E3QT0yXPj1/lHFKkEZLsgsoZ3a/K3lkYZ0+sNOa
C/xY0AaCz5yGA54FENMxoMASQq1CVs0ogwy1zW6WxHZ/J1BmeCLAFzPsaqRPnrDjRpADTyjzqZUy
G29aDsrbcZH51/SlCGNWoc//HzHJ1P987ClFxEniuzR3QxJ3uClPdwU4BhR5H/A2nc1p8UK5u+iT
qaIcyVaDyHn+gCPloeNk8hBGbyshHJOYstq4YeY+PD/UThwTVe6cC0wfHI8zizy655wqUkGbic0A
vSzLD8hwjzYU/jXtSSPjexzU0Kl9bYZtuSMgF1cEU01d+8fnjEzzQFXZw/XdgzBEXtnOKfXVGwO6
n+Q5xHvIJ7Q3mzpXj0yVufSeDlipnROszzgPbnQsgebUUoCVK/vxxfZsQ5N3yb/ZJ3Uhc6mZCI2k
pFkAOZSjDxAgq9/vnyWPEuWThf7W1MKXhLEW0GrveAYIU5epvfPTqRukmOGI4tUuzYo1T26O4EFU
oSDRPz71rGYUNP+3L12nlufjxzvKFmdzHqBmHOQEWoRPqVr5uAIqqjY0XBu6qt+tShe8QW1UpWTy
N6XDt8P4pRA7kEgKH72v9vLKa5cC+2afZmT6qzr3PDqJ4Y/H7SHwaw9RzPXL2QoEEy/ijmKLXU+Q
SE+jmN7WThHaVUc9Ls++ZyZOnhengQtWGdhTevIbLGyr58HJGR1Ka7GHDAZQtAkygdD7JUPOZwYL
yDpspdrij8+IIOgCFoWgMKMeko5VmX2xEFV74b4S+HCQ8Qa1m8QYvoLmBg5NQjUHtxKfZpSJ8tFn
OX2TGE+ZR1dkPdS4WtiEkA2XpFNRlzZAClQN3Nck0sSPCxxBsdU2bWphW9EKAh05+EbBcgDV8Tws
kpF17z/UlHBEVgXYRMLR8kldTyeVmT97QOSQ1xYB2p3wfSEagzv/ijxORqgb01BPFN7rkRspPt97
XteG7s2v1I0DJnXituCCRbpt5ZxicQHClXWfGHUh5g4q7Uf3Lm7REJdr5hCLKZRweH5LIdGqzHvg
mem8i+IhHKGaxFaVHZBcQBTfFfPeUcQsYRLWe5XWTPHuNM2uC9CzWktjI7jeiJwOOAeWgF8H9Rfm
yq95Gz1vHfMgKMJKhJ3IYkXDEAG3Cso28wXgs+S/fsWWnVaCvd4LJjblvMq3YH5jreEJ8wiAUOPl
TxWAce0moRxXT5aafoyNhPBVXltdjgL6XD1McyYl5leA2YhyczoOPZC8br5BaGM/Fn2yUTuaAJvY
kgyoeZWobTlQmzKpaweQs5mUiXkJDqD7rZsICa//h17oJashDgTlB+2iPkFO0CkOyUTvGyQocn//
1tkLh4hlGQvcmLIZ9gqN3sheBUhaKk1J0xYRKZ/itPzISBTp69zQHcI83izaiXJELAGsR59PqwJ+
Yn7yOuhTlQIrM5Y16HcIRofwLVOTTxzV2AlZ9Bv0FFNKVxzPWmJBtETmG6LyhBnwiL0Ep+7wqXgA
uj9vHQwGKAzZZL7sDIkCgGq9EnGgQwo5emGyYMOrUNWUgr2aMma039dDuoqv9b4AZeMKJTLyNUv4
h7XeHT2Ar/7v0B2oCnBKXSsMAE6d4R+NXDL3Qh8imZh+bCgjJwn/c4O17CUdL6PwhpRQEvz7WiJr
qtG+RWb3XtdXEFDTlvTt1VGEaACZlb7ykC9b7lOR1CcLzJApd0I1+euSONjLreS9dpQDb+2nKowx
56s5Vg/gyeiylIjY9fOkW29P5cwdCraikNmvR306EXLyiufaHcOt6GrqNdafp0oRYLxBYve43rzi
+cX/3LYKJnPAKZ9gqzJItLsHHW/PjjjTsqX7PiYskuYwX/AqIlvH3cqGP1OPxkkV67JIFW4QBoNK
Yn4ddrX7c9uCOwZg+CT/9mBhk2bxQYPWIDT1Os12N62Q93m5rAfKiz2IvpvLv24uJy7cIv7tBIeN
NSi4DucO0v3SHxNFelsIcvX7RgDY68muF41UX3qhASCsMKck36lfDqv8SzkkUfe+gPcPeErOBaXn
EV9is4GGgcI72m8Nu0XIb5gkOBWpHMmNs2fvPIVgP2p9PEkqZr7a25Gi772jxFGItUpdestacA9k
iRgW2cQ/IPyn920RUUsR9CulwHcChO3OV6xPzlasR4ffqMFCzUvF1PBWW5TY8QuKnq0qdF9Ubhen
oHZWLfKcCdWPjamvzV213G7cKAFD1Fbm08LSQZx0XlpstR4WNxSmRQiZQ36ek0BYuyIoJ7oQw3az
2O6wM8+QPJST0JlsCmPJzK1bg7Q1vl+yqzHGy/Mom+nuQe1rr63Sy9dgPlfxkjcDmE5WYVc0SQVU
GFbpsIQemPApt7SaPBUSZLtpDzYJYnnPucsEMtWlfseOTSlA2jgrHAdI8T5YJ1Rgj8eLbH2l31N8
wXVwZpzf8J4FgbheYVrT+mRPA0za+qTiz30sxuisy2SsBLzR7daNVljNhefziRf+dePjjGpFgY9+
9w4wmAXTDzoNrlwGeVJyrPjnLlR6EQA8Wj00E3bNKbHBlKpj2Et2BfW4xQJifrJ/s8ME8nOG85hk
+Ov8g+ZQTiRUlEc9zAuxdQUzycnkfS8iTFhmEj/g7Ayrlx9VZNbA/ZizotieJivYUf2Cva7KemB6
bE2ISetKHJehUn10b520NgmeWuaWfmyJjdPSoLsgTbBJheHqbXLwodY2ch33DlI7by1yiU+OlUjO
3KYbznAmEnsUQg2YlZgPID+NXfHTQcFDmhezdRrZ9FeW5aY6EWWHVzF9s7W8KQgRUJy3O5Nl9MaT
Ti3CKYU/juyVaffvUW2hLRzChv8Aul7zLu5k+0rc9vaBL3JEvMcyiR9lKE0zOU8QSM1DYYJ885dJ
k04Lei09CFklA3yEmU17amIegcAsE19JdH4FofFgb9tgX+zAP0KHeaipm9TxaKSDmNUksgNjeCaj
gFeIdfIIeSoUWgIWLK3spRPzAP9p4D8ycHPge3Bt/gFiKyaTlbUwXsCt5FowaRgVjNwtoD4zuJMW
0iOD1Mxf1vomkIZmRaW7NReiqDdvOoiSLicaXFDr8wDPRrHSXAFMnqHUsBwPLvw+ZAOMJD/PHPSF
gCFjlupFM7uVxzxBctGb6wEvdsjVrw9zjUWOZLM4PdSOzYsiadP4J2R3HWuhJdKQ4oka0AxtmZJd
Q8SW8SPR1Jl2H7c/3lobmboN4E6ECDvTwDkJt+HaX8Q2Gx+v7mCNYKIGLtRE00JlW9kBR3T6Adgr
yS03ho8hMufeuN8AZGyfqBrFIU/P7MwG678GZLmbEN6nbFohDF0WFLSAJG4yYAPtbunUEyunDbBX
tsxK+GPLJiHGMcar/OJ0Fp/I7+q5AN7IX7OFd+ZBdkYih3pXMAqFQvOA0IInp8aHWmj5I0auhHgM
IQevH21zIT55K/aPBLW5eqCpxzAIkkdAXeGISs7/Df7UKIg66ETUkiNF5jhJ6/QN0L6JFyZYbUgp
KGA0awepX9rAyZ19RB2aPEJl3OcJrEbuloATkMxf7upu5Vrx9NuRBP29yvlB0eXDOMXNPquJ0V/A
bcBaWdyl+DDB/X9evQ5n4AzxRNSowcZZzYmY9WdUfYHfiHOIFs7aIhWagNT2rhbvu6VrPa4PMsyL
ugXb0rFvBmLx4/phLy3SahbwfhadnP3PVcOH9GvvVEi92wWHTzslDuDe2JEZEBv8Ei2nh/A1U9vl
P21KW3vBKE7upUJx5u/OqxirVRIJ3LH2ricewIoBmoDPNl9Wd+PZVXDdqy7vRbiFB7g7Kvcjd1Ak
zInTwX5ab4OWqrjjdhu4dxLwsvXq550AElNuXLZpIueArNqq4is5ZoAfu4NPJNMQCNihx04FsD7q
L3JINC+kanf2nkayNaA7VTl9dpmq1i5sViNv9s6gskw6yE8rESl+AQILUJj5L/Pf+yXpElPTEW4n
vw0sN37AJq0dgvGrbgE37cq5L0LvxHHkW5Buzu1thAb1JrkbWEcHBdcaEMCxbrLmv6va11BTwTQ6
PuRv6bGlAzzPp9O4yJeozIIYmIbJXY0yw5o8+M/tGHbFK+kiq3B6FbNm1fRgkpy+MZ1ssE0UBvS9
cCSk1tc26H4OwFa0vIIIje9m1z0FOVgSG8LJXJG90BrviodTG/bKonlS/j/T/Tj+sxUtAldstYZP
pDENW4A517zk9cGZRcwOFwZIcytCKGGzG8jU//CouwEnPulbdqHI9ypoUKcfxhumFh8EsU5IFmTV
IwBzV3MY/wO7rvVVXVuO0/uD3D6PvOSN6djygyVEAAuouxhQmtzJO6wxeWW+M1Tl6oBGEYEzrp+i
XkgYcXgnHkgOkrF9gtzQhlhRJ29CYuxbfV7i3c1WZ19K7Bnm7p9FwhpZ6XQ4wp5skxYjAmkzRbT4
lTaJtjiWTvslxQg+0Hk5jdYmKuNioFNIwrPsGfdM4bs5vnWS1G7m/SKDXxeK9hM5tS2jl0+gQEK9
nWLGjvb7ccfF2gq7zgfDaA1091X7PJYnY+jZqTevKP6YEXLKzIvwqhpNfXKoPRQQ/L7qMlQkV1vW
5OfBC/PoGiEj5dhVDvFyYynj9T86nkzZUX8meHOSLbc6Sy1TdmTD6snmwKAuC3UDLIYI7IneWW1S
+p4cR4joz/ZeqZTUagSc1lfI0yL5BACZcrGxCrIkN1WW493QkzyorKQXg/wSv/OtFfw4BxtOdkio
64Gys91gihMEdi0abnm9sSxU/QpUHkdhjUChSiJrB9ekjQByTnVV1heCPm5TkSuAtkpZVRBwMhPL
A29GOGsnK/1xv8gdJlddDNBd4qYpLTyncj5sDtme7eeIxRpzELHyIkhBOiktpyrlu3s/cs7C3wOx
sF1XfxSbmmdOPAzTePgemBBMxTtgj8f4Y9LoNmDN8Vf6NaDejjHiyrl+U3p7PbH4608pXLVJuBvZ
s2fymos75s7gvVnPLyGPpL2wauVDRnmhNVbH19/rOlAij9LrTjRXkaYQxz34RM0rTkKQ/NaelXe6
nqcyw9oFtVbDELW9IABZLTUApSi/gynETT2woql8GxbMlxA9uGTFYa56ARCWmAqQ//dkMp33+g57
CkBwT+iTT8m5WWed1NNkMeC8AD3KkIPib4FZsZ/ZZn+npleDtdzmWaqxycl2MJwuIWtQAA6PftDI
a+swft+ck6ZMYUFm8hgfU1ovoe+y4URFdGvs2R78vW4mho7u8j5tAtk8oM/COdzQgTSDFFtQ3mix
zS/XEegLz2UXeGZGdD4g5ML5i3NilgFA/Vnih0M5j9SVcwmDHfXp8jy2JC7LpsblsS6D3uCQmgQj
SbE08L6mCIHwsAAuj1lfMVcOV1kJUJ+bV3y82XYWazILntP29TZo0i18nzWVA1CJk2KWMTIWwKKd
j1nhcmUjj9XTosDXkpsEeNOPEiXD4p6oIaejsCW/a4rB+Bhe5BL5G7W2LIKuihIIuzN5CZ66qaAB
HJ8GuGIirUNtWzywOZ1m0RpbYrC4rgvseBLknVHDklyN4vdvklEIHLxiVTDOm2iwOaetx2y/FNCi
ofWogU6blSHlpKNfHC9UGf3tiYvtRKFACNXYKnRq19+I7ysLXV+zUHT6tor+n5aX8cMhFRkoN5xQ
F+qUEmFWwlgyztCoGue3Ykn2w7Hc91JArb7aWkUggtHZ27jm5Ll0huj1QAEafsPjBs5G4T1D2SNz
ZH2Qid4SD48MPkYVhHu0DRRn0UJvZjgA3wp0Dh/8zgGCZKnMD5UJib1mLJKx6s650/k0KKA/tQxs
EZfULJBCr6lk0x7zPgpLE6DVg2PyEYpV+NDsqNpAkB9eh1fg2jsdrAUcINNZfmjuz16lLxsrMat1
yWt2aQ6Mea/aJMBOrmchL262JkiPoouQ+o3GFUEF+SAMyQk1AHN5ZKopMwsp6MVJrT1l0GJsRvBf
385G/miaVeWmOs1wEg5qjOtc+tnqxfGscVkVIYCpkT3u8PweeD0riW3Z9aqqWnr3vbsX1m+GbBG8
VSyDCGeG0lY9nHXJpsU6npZ3w8csnuFYWKJt7pnbUeY9oPmT9COosbBIDOrNRVXGxaz52HWkxgCr
EvGOijdtWwfCKf6Fd76OTOoTDd64VEdgMkAM2nQ42gnQ1igf7ZyvIDZdgef2VLm+OnMOpLLtkF+Q
kiU8P8YL4MTTQ7w/pyn7jiO/GcsA0TKsCxsx7ZMYUNceL1UELHJmpaV6zOOQidpJ+/C47gvuJdNL
A/QYVdKcZCTEDtS+vjJR93Lhb7cughA6VWOJEq/eodLMp35uZbfmiGZXllX1SaGx9DVGNX8kjTNX
r3elCJ8X7gueN8JpLv6c486Z5H+zaRVOb/HelD9Ndx4MIFwey5PN2B5p2DC3+phDqndPmsRx8mN9
mAYDHIbopf20VBuCma6V7VWArwWgQHG5xpNelIVYaa7bdyxGHqcXYpDR0gOBi1hlK5hZluIJQ12G
4tEjB6MEzE4FRcBR0LTKr6Ks4KtyZkqC+i59LUejN/9FST56Dkit7LnFq/29NRhbYFwle0nkku5R
GD9OGu/3JbC+LLX7IgpGx8KHiGoRfWjc04Pkh65F1MWa6s1+B4ov4QNtBnzOuSg2ytw1hY43EVEi
yr9mtqaqdE4nGQpCfdAQM4S8ZOGeB7h2rKCsK2S0pUEJrPAeRUqMbEC3dUAGcdNK5Wo32o0hKsGF
GfOAJjNQP5jDxexTtqYQD6nF8Jd6v342f78THhrW3XHBlH4/3iNMHSfUTK97zU6Ix09U9BCIfTs4
5FWJTr5FvbufHzV7QI6wIkRTj5TIw0hE7WbP9rOLRom1+ULNLrd65fIwsOnWXieyLscGlyskLvhV
uKUVPUlrDT5heV3mTXmGUzQbGGV+qsEEozAHWt9s5BcC8IYq1sWU9B8CheHUzwuSWsWGjuMWZLcx
Ebpy37hAXsrq+KSjwci4aukW32xpY9gFH8E6YC20sNkTh9R3VlxCdTkmtfuin9nmFyHuZ6ZnguPy
c4+u/VK/xYqlE3bIIDu748IoKpslAb7k4asBo6b0FthCSP4TwdWnaVuFonMbkV+uNteu5yni8chC
ShfC7enSExSyGcjnfV+9Mgx089BiwzoVLf08XqTHtJT8y8FsrdCPbgtlekyodkxdAYpJ8kmaQGel
Fxrgy6NBPT8lNw/jZcOULi1gdzvWk+hWVbHjv/vs3U+hSU30ylOEsyIPL76TsLFGNhBpcgQ7O+mX
kDj7eAs0MXMwHEeXV20LxmgM0xDFs13As8v2xY5Ev34vhqUqMqa0W3BSAWqKbde3MNw73pufBmke
9O7kFzHbRW3sPNvqeSvSej976ClZKE7ZBEWrmAnU3ZgXkXvY8d6tt64TNfYk4hH97Xtn9LNcoYE6
3CUxTn8cU6gTQam9ZvPOE09rt1bTwZKSeParK5gvRvG0TbXRgXng8Bh/Tnf497cLjBnBQiSUGvS2
htDT5DoUSKiw6Ktrv/sJUg8chqLJuncwqeVEcTX23tS51yvZO5FQ1Fuzc4GKk/BQQnOXi+CJnxEH
W2+jHw3s6qyB0FC3aWESk2QjiODsR8yPlwDk0i5hxjAyMPKW4ZvFJKONS/RlpCrfV4cpkXAItq/f
HGJsJW8mrbWaIrKHaciiAeBPRQlkWfLDedk1ZDPMxT7lkb0KooaXlQzV9nv2wqQx2IPfB5arO6VF
nKYQjG1lH9wZ3EefjL56EDv5JkJxstr61jMvEMKDq+7SdgDOKB0kYf7mbDMRwVtTENT+4nUxKwhD
dxodNJXrcjo2V5hvPwmCeVJOdnfOdeElsvKOD8l13A9WE2YlYHlW4g1ETKrCEhtm5WJZyIDgiQ+u
p1PgQN1xmjib4gtrIIu+tPJ646sD+eJmKOa5ehgps6a7pzkvaREa2a8lvbG9BRBxFgB4j9x/HKVy
RpBDP3150fvJafYQNEbuW9bwUpBcRQsJpK3OpLpSll8vn3efbufwtAngMLpusisqyawdzYrdzTPo
Zs8USk57FEXPH/M0i3DQsmNJ/fpi64kI3Mw5524kn5hE7h4vph/sEgumjtIM0iKrPnTKmCZbTZzB
FBrtsZFEPn6XuVRozydBDbIpOb0SSvpztB35Tf9h240/u185wAzKVH8pZ+IoATck0NVYb+1YWBpx
/8e72RD5SH646lnlPX14aATGdt+g4fZiWGnv+1yNBKKCaDgWua4bNpUyqB31ert2BMY4c+GKwkU5
Yx1F+Lu1EjdpbDsNto2kwycCTmrcsepvBrS433vfJ0p+Q32AHeIlmfz+E0Z6H+Zxr4LXvz+eaGRf
THRwo4rzympzSDH/IMhmDveJrsnDiwr6eU95HUwFHTyH62SQOvEWeOmDCQrkInAVhaN59B5oo+tr
VTBViWIHxlGVApAjKhWNaIqrHQJz/kvrfneekD34lr04H+pgqHVBBG0wLcYu9CReNhDgsvzIIzoR
nPThuHpzWP2powJdqCLbwYidZgu+mUyzRBQ/ZHdZkRNW1bpSC7mxz4u1NnPs6e0NaXP5osEV3TgW
8Lbsq7TYHa9fA2c8xyz7j1poPl8wXh75Scl8F3QMv2jaIJpB3rlGceDSwy+AXe7s6aVkAoO3VUb2
Hh3WGANbSbF+adXOFEa11+b08VvwPwGqqXnz/eBz2/E+RTssry2mTs8aG+qkX5aUPlYdc8i5TAzW
msh4wUmAM2q2b30PffItb0SR+tjt32KohUMeInU1BwRjWem1zqYlGYDYPARhn89jmr2cViO2A5w7
8VNJ45zTS5TTThbievISYmacpG8bFOByALO5z0yVPOgvUml42lzweN36LR7/WJzcxFbyNKVDO3kA
UbiUPdafMDLUEMsR7YnMtP0C3TIsxIygvsTo9pouf7UOUfBu8d+lVzYi/8af9k52NSJtJPa71+Bq
QTEfN+vyTk8Zp2a6ELVN5ikuYaZ5qZtQ7X8rrJhjWgonrQ9oymo0fK84eOpXz8gbvTLqF1Ql81p6
7mGJCZFBQO9sH5WnQla08YPjWRJ1TG0Iuv76T+NUPmOAK2vU81UJyEynUJDQ2DO+bXnsR/YkTY4v
4d8oV0qb1vdFoUrFixxhKP2UiGUE58S/xtg/gGjE+5mkNsZWc1wV2X43y1tiaNUJLDN2m+FDeamT
/krFKjlWLi1MMYB2ZXdGBcPLurzUE3vhQt30Pi7ONoYok9DNhgLbMwO8Vf4+6uv3Ie/mVjIEY1GU
yeuZBBxh+d6ItLvUsqBL7Hf4NZ3WVbQlJHvdcggRway3cJM8y3PsVymEHWcL0zzIAXoxX4o+g86n
GbJpLlvZ++hHqDwqeFDrgGo7psZEod64jQsH4kTg5K50WqXaVpq1raFIk/PAsJdL7Im7zNUYyNjo
ScG3FywbVvNAkdDg+ESV7OF1vzlV8JL2VfK2qRqLGbGe+cMRLuDaq7kXNlaw/02sEH76JidfvMGG
nMk30CBycuALGCZbUrpGYL/BfHVmJj/WkbMpQ2XVHp/HeypPP/ZRrzXQ56uIG0UliKTu9oddOeg8
oUZf1KujBLXDgZdoRDPLU7IzED0SG0TMMfPjQnQkSei/DMw2SlnuNTFFM7SRufl+JifsXuje8SWV
AHKCRDtq5vLeGQ12mel0za+aQvVFPqKIaStqj85ujRGKnn7ovhZNZVTRMEwuebfD3uVnw8sVRGuP
UXKZsQZGmkbWajF6z8QQFxbUcBpMkdc+PSOohLPumBCFA45ZXVfPUvlg/lzge6xmWoUBjsqbT512
MNAooB1rp32d+rGdwicfaSLvrYi3HMNF9F0WARGbapN6T169OUiWc6983Nf26CyrtaZjdI4nkIRb
rhs7J/Zo5EaF1f4JzfTSo3iiL92PInXf59zvH8zB9rllr6h/pDB6NZURAxBxOmrXBp9Hy48FZMog
UYtvYJwV6u7Dz4nt5U1cegSKVVoRuHOJogt+uwXVdsqHYljAVvDhiw3a1ehc6QWcrSzeIZtjLgOe
p6vHpKLSQTgYDFar9/sfIqbeb15HUfrTQCggeNIXQXUu73hkc/4DHMUHQ2gRdEW5tJIbnd34M68O
bK0g7uEKdjgNCGgryoID8Fp9rZjht0Bx51/o+wrgGBXdPo4raubfRt7yJEFkx9fhBUDCwLos1AjX
VbvjpHqZnTAUCzK3f5PPE8af2Lbh3Y2D600RLVhbw15mfmnt+tLhFUGoJl6MI4JLVueX+HMsvBbQ
KmtaNtdcorVwnTAlV4nP4ZM8DCXrQUg/ClmWu6gberOVp1MgRupNnuy6VGSaASHPQe29cPRvck1W
WYg/MIgA2MoDSGVJqlW9bRVNZeyPzmzWRzWyRwSVTdbP0zZBt5eUBdEVQMyfQ+B5D/l/siQanZKE
PVfyXkplGrUFPHOlHuDpfRb83ho6kS9bCy8aw19j4j8xMY7aqptTRQXHccMAQD2m5jT0s+w5pdTm
+eyhjTm6JIhy0Y0KHgXJu2tU6yRgvvG60fkKRhtyF7ChTKBWxZmd1VnaOtkeTm3IYQdQUdni9MjI
7ThGILrBL6TwAtydhCNYFlbXKkMlzFsd1UMcvhXil5JwRtJ1LqjPikL6PScX2n3JJqiOtvMlRV0C
Ru429NoxpZ64rLRgaOnuKVE7PF3rQRtzjEK3OuHCHGqvGC0a3EEYF0AKChOMcrpzJvCfS1UfWtz1
JhL72Q8NhAf8q5wZ0rloaPzID4ioN9Pu1Ad6Glm0gztS9kgStTs9MB/GWdPJMgjk4DmyVKyaheE4
iG+shHUSXlbQjqIwaj0FmufhxlSIzJUQNCB73izthXqQLhNuJ5RV6a4b6JqiIIarR2fuZHVr1Y7C
wWrfivh+aN41OtP10G7QvqADOVWPrjPguzSX0PjtPowOWTyIQZZUptNR+dK6s0hNGFjOl0Ddz2Xc
7ZlBV88EM5qbyQqbR/8omVtRZEw4X3m8bqXop6E9kcJUuVbKXRJOVL3yNJxckEoon3PjWFzgN+ON
KCZH3JEcIrqQ4UqfDQuDthGpvvk9lnP08p8duK6WWn0yRVbvgdvqIQH5mqDyj/dkjUB1HGKPFwo7
7MVFosyfeUo5bO+nxPgvDF1PrHIGmGhgsZThWBK/1NttrqaFmEXZrHOSz6mC/g1bPg8RNnvYdLbp
qjGhxebbGFr9i0d798X9o4RdHi+gP3I9vaa16HnbHkAzd01io3CN2elojgnTT7ZR0KOsup4p1zWP
4eDTmXHTLJgJV/FTqzcmKl4YoUkzvFbrSsKNI4XhG2J+ih3ypKHPE2ADaI6KL64Z8DlSCGJCrI15
nKxZZ/Hi2S0+ox6YK58EpzRvXy1WG3i4h4aRBsH7rvPBFw5MJ3eKuewFrNG7hyvXHqdYib5sh8S3
3CtSAtjmWLcsf6GKUqBgHDD3XsBq7ssPgb04xfb3BjnQCTVv87G4gc5KQ9VBsxllfvprA7IzpP2/
1Z4fFsKBmoOTIJg2fqfTJpfZ1MdFD8ZlEW5WQQUwG01tDHiokFP8+lEUSR4LGTA4BviGCU3B2u9V
nmfA3PReJRJLlVsw3Fe56awEDRkEkIT2kPb5nmnQWsutWHWcqJd8fOQEtq4SGTyQ/EFT7fao7LAu
CnQfZopldak1ABlB5fXsWf3rE43+ajQmRuzvUQWO/hkUdbvo11jJbFA1K7e/qR5hELOJvRbIm0bd
3wtaTDMmd97meBP9ZTbgTXdVVUCpzt7TGIMLFfS5k6SDgTJwetjtxQRqgLU9Ie/giyPGQZu/NrHg
G1lrjt2mvPWhR9M2AIqSvU6El1w6D5rliTp0NvRF+pv/c6MQS8OO+0pf91YqslXdMchr042WURph
XAbnhFhYO0MyKjRqI0erSoWMZWPMR9UhFlJyfbYpGQwutMOGR3uvBGiKd7zHMmiYpZoUubCnIef0
7Xq22fZAwz6o8kgUqe+aCR0edl7JPax5ygQ90A5b0aLbggCvajPBcEG6QoONOqUhBAbFeyHTeFkl
CSfhjowc+hZC/vG+bwFKOfP1nUYLbjosV4295/LWnJScR/+R0DWwabIee5gzMZZd0ISfpBw6BjU+
MwdMF5h7WjADRtpcsZzU3PRUpi8IZRjnOD6oSqNaxQqWy9kifzuzfCQpNbvXVa1VVRI5y3QW+7/R
bWeMXbJQQzVU4imXPxY8aP9E2P6MQI3rMPGD3QpRGxfZoD2/DgOIIb0F2DzQgxZNdGjDFLBOA6PC
a4UlMrP5QGvKHbraV6iS/D97+cSpcTPAF8daDqNVyDIdpwZfuPQO8zBMifsXylWomRUzYpC0gsYL
TzsBee5TXNDJRaAtfC3h4+e+kRiqnESTt+46yWVXIS6uvtlmqV3NyFSGtoQL2zDkgJ/1Jk2BqAkJ
vAnu+i8QJTF3QWbhT0qebjnb8sY/TYIgIfQt7AOkabjaGNqOjEJ3mgzORunIGLKIbtGBJD3d8hDq
vYs5J8CGqOUgJWS7E/T5VBPohHR4OfsmhwOeSxJ/rDqnSOIGk/2nYy2KVwCZAfrmGeCX56lwxyVx
0MYlkpqUX7CfJ5LbdI7T4ocol5dYpMTc40OBJwKKH3xi2KHn5EBUopw/+1mWBvmK6YwohAR30KgX
p95CdC+OgXtmzMFmFQPKjEUuRIFasc0JzBYqiZ+EqzWKmv/yL4JuCJnz6Q/lHamG9Ogo1CaM2prf
f/bAIkzolZ96voMIxExpAbZNfk8sElq/GJBwaxgWLuNLWojKfTvsRkQ+KdKGOuNIHLZXMqOThbwc
CkPoE536bdkg4221wv3e/KPg3A2uZKkoeMxufBMFp9tFjLwG5KXFh9ghB7uEGabNbkClzkadj/Pu
EY8JzY/AjwuYl7BZvx34YtNkKZT/5neYSgno6T72/AWgBxnQuDk/3SEheyutCytoLfBth5ngHIeK
wN3VTND/IcgJUC8pJoqW/Q79k8CW1qKjT3qqxC1z1Sda34PJ43ggTrG5GnT7nreWmMmncwmlp76h
2bG1Rfgv+jpcaAGMo9tXOhUx6qua0H9GG1eldmecIvhO3F4I0vJ1DyyxWudc+sWQJ7+gumng4dVi
o6bJCgl6PnFTvlnB/8waov/g5Bxqhunue2ZmTnRrhUQo8y3z5+fNG2ayscS/tU98vCN2B1PXcmpO
rFkpCMluBR6Z2i3nUXVrVGaf9UtjUIIK3xZJNJxphhtqnqYN3mlVuSdoUq3lPTnC/7/RUK4Iy70c
JJ4Fbfgm7qeU4BsLqCf2kuvap55V8mWE2EAZGhgvazLznGTi93gvHIVW7q2UVdZgJTe8Cgok5uP7
BS3KGPBoG4XOBq6LUsm1CDahacspGXblRnEfkrl4ipF/pxvC1bzZcR261bFOMdmeac5KDeZxl6cf
gbBwgnGsos1QC2YS3P96Uc4KfLUyG3lZvoxRckN70B/FomLpx0gyL8LuF5LxQ1JxcDnFmTBG7E7H
lMV9//hMZZ+uz103d+RqKfdqeBZqJ3nrC67ao6uNRKuIk1mYUxbTPzjkz1VBskoeMa6kCn8VRAsu
IUxGy6pFvqs1ukf5uKv1eu852Rn+WlN+2uvD+IGWrmVp5TIzsOGcUPJ0EG9/sKFJvvSHay5f8yck
LOzeS3LNYW6meDiJQ5N1MOmaq70et/5JrrSz3b9H/SjXXLLcjSvOGvldD/aw9fXNbvyXYNBZt815
ukbzziySJFJmax5G1vNfHYUtf8nYNsY5gyCR/pXh97C8B8LUshuBPErK9+MOuDOwixf9CZlkJH3b
TMqbQsWWhvRst3kPzdi8kaW1BiW9FXxr4DvREH5j9kA+W+RVhj4TNrzc1INWB2ykmGPihpkoqqgd
kNCpR08qjzr2Ia8I8jayM/tuMtFB+kR0edakfwRh3ChVWOy1G07P4atlmEfTyMMSAH53tuRFo/2I
ngEmf6M9QWSG46v/GwffpO1DzJ7uNOIEZ4oA3mProE+CmzVHVLASBmE1RoNvf9j4KWr5+p2WuVpB
o//dXaPywrgJTduM3u2ZB58Ut1Q+DSkfUH/RuevetUAvUTYlStUKFAd109HPvuzOF99vRKlO1Xgk
VYZmVVltIskL0552zDzcYJDiNICoLfmUlGS6jzCuBhHVxqqTZJfL3jo3ROBVjSBW/o+Wk+O1LY7m
peNpL72AklABRN6bKx6EFETktX4hO7n7PmQUWtKFgBVplcBKVGLd3CZ2WbIVtgCmFkB2+jLev/U+
0DYWrGeJzQX1fgeiaFn71bNtlSy2byuCHEYNHyzvA8c57DMrWjPF4z5uY7o6VvfUbT/sDd4GdWMe
xGXYhv/ifYa16fyjPO2SU6J9r9wgpMhFTaX1W9RfqS/kDHdDPCQ6L5Pui6JGsF7WEUym/C3c0wLq
Ap7urgIc2Fn+ceAqd2LfkIEnBIMs41kr8WbMyNqI5QNQOtsoJdBuNYrBbKLxu17dIpyJJ+oCcemM
PUIzs/wJDThINCY876onK59b34NSFNycVBBeC+PMrwkqoWxpCIaHnNZDMNlg5wQVvHxupO/X0z1a
ksNv/wGMt7IWvYtgnL82MyPOkV369asDwtOVwHI3JcsFt617NalHkT4KqL2mgFTFlEHOdMBYAZ7L
ldC5q66qSkKV7BK5WlwINi1NjYkVoFOy23c//ktC92BZGqhFh4e+6ZNdjfuqgKsWtlLkEzBI22bZ
8MMaedzdyrBTRyBSb2ObJqzsJ7W4gNAO6UIfxUXOOuRdPy6e+WFbMKamxD7R6qd2b42dZ4zxvlDt
mS/gMuiesiXx57u9ZAeRbPTyultpZkw83Obmj20my/o503SCoukYEEvKLOWmF4+fYt9wU0xV1N0V
aC/xVJfyXzC34/iD/khhGz0YgmB1mtYP8BcP69RUfKzH2MdebT14MxougDwvBAiaOXb5uvE3zLa8
gEWwj/iYuznP1GsUC5RtgIygYPY9lNIelA9fLeB6qUkp2QUclHlChXQRm/iLTZhMa/l+JmJGuyI9
gqx54G5VJy1MOzVmfn2cZR0EyH0TBZag0nxpP2tk0JoBxvC/Wmkc5GoUH/9foBlWTthObjcQLSR1
/GKPlAbZHJqcMVxdptiJdnaQfnKFcYcCarVjiu1zVrb08ytyvccs+CTOyDAkRc+Vv0HhzkTOxhy3
iQxsIuyCFXJbgSZewQa702qVbOosFRsHsEuOoJYTLdcO+RLISpERyaOJWBFb113noYe8WZAJqNGB
/bDjPYQPNhGadOK18ZQtiA1RpBF5i0ONQ29Z4ADzI6AeWMbqXSoMYmuvHub/6i5kRrm6FfX48wVT
PTojNiDvw96UgIHRYN83ZUBrgLhXFV6vA6hrcoraHcxOuFS4vPdWxWzxb2lBbpzFsZpzEhE6+m9a
LkOyUM6hNyAiq/var/SMgTbxElMLzOApv5DgwDCmsTvqgh3LtAOBpk/a92PdbCZdqP5JbWCbKpJe
gtOcg11viAmSR/jbYotajTwFv+J5yzSa4R58QenvzISw3X9e8alonzB1Zw0fu91mHLWcEwfNgGGv
6NlWBDcG67uKec5vitXeCQ1GgTAgAmMoHrIF1u6hyYGuuQjCsb/hVuHUGZpJTDx0zf7DJvPm0sl7
dDVPn3vERVISgOavUYnsm3IAXCCshtXWkbjknbSTZ7b0LV9X0bDkrtyydUU51M675T97cCqFsd89
Y7Vhiw+QzuMROBF6OjbgGsg77ms4CD4COr4QY06iHZj4BTDfXEE+ks3EM7/pZIkBAC8cZS0wZwxw
vEipPZLEQzgG8lELPfuM8gI7dEH4H5fsljFCJy4DuAkt+AMoqAN3wH24eJLj2hPpmmyW4UU0ixRo
ekCvug23SlUt5kMjr2ffP+YxGZe9nR19SZGXqgWhdEvqIjXT10lqLDdwIthp+vGvLxJMeIlTKQQn
uJT3ReiXPKq60WFxfk+5kgs7a8OU/+c8MLzLOVk6uZRjzJZvt39L2n0S1cLPPkQgMUtOQjOUpm8D
bfvTSTQsEd+4FT4CyYCTf09x3kYZc8dGevaeOdlXcYMcDB6eXrwto7Ls3m5IkJqKD76omJaGWIOb
ZRGpCXuLtn4hdqUhaGT8Vg6FmzzJe87e8/r4+xiKIyucJqqojFxIN36fMhAH6V7sCpImREzFTwPh
guiuOq7sAII5RiofuYZoSQ/IjXczeN2wpTQeLWSDDTrYzTanYzKMnSHTBx4W65qhWp8rHVexky7Z
XzlQygNa6YnXROsok2H7psj0Lgaq5GtlnNf1rBs6i2cSsFE1OjRlf1LasVfVfwMFrGrl/wVX4e0/
Yeq+iAonE8MVASCP3LbfG4fGRdqq9T0ECNj4yomxrsOpLyVQaXm5lz6NzidoNf+fZyOfKf1v/bWU
rv0srlaC9QFIPLoUJTDCQmARB/LAP+2k27f5E+3OsCmvq+ICGq84Vaxh13NbGEIXlXCHQh/qBq8F
hR23Ul+hDJpHLNmKYb/uKLJzMNPSldqnUOP7Qu8bBIsMajpH1IaU/CJ7TlavcUrxGznCa6ozvkq1
QhPqFDTVT3EDzN2a9jQ9fFeuifqPiy7dmiWOK4OZGjxVze8zrN5b5C73Llie+KfTZrVbc+aCz0Bx
OIfKBvR+Iv1u6vxrgpPcWF4t0eUZu9Dt/6Heft+7yZ8Vqp41MObZaisSepWV7YRdUXoAC1n85///
2TQYsNZ157V9rLrk1rH6R+giXCsIbHcT+lyJzPSibOTe+i4RgeLGUB0Qbs1sJXmcfujhpHKbZppg
l6quePKO+BwvZoUhE8+zSn2LLsryNx29XDxlancChosZDJdDdeUI7YdF8UZoo2ZlNk3sP3IiumFw
6HjFgiHiupIkAt1wxgUwM8ZlogypNUOJzjbyOqf9Fw8Sz3ZI9Bxoul5YavclyMArEfPyOnWiW8Wz
OTQXjE1NVzIfM6OcrqcZYRio1xOWda8MiXaQR6+QacEBR0Zg8+a/7aofwnsXEPZaJxCDIiouGG6F
kv1nx/KtQlIx6eRiJKAbHxdOQfJH2W0EqJvLFJR+auM7IdiPDMPf0iUhV6vei20Lx6gRMroQ5pRz
PiOPk/yhzOoS4gxofNvzFYptw+wHpZVus8fztw4BAsLmsFzgveoecucDAFTRyHOXCeyocQ2m50j9
/Gk1OxCtiwHDkBRTlc+9V0AwTevuQWUcSSToWQaZ0UfFx1PK5lIH0nTRI/dSoRP02i1DTulJX/pJ
MI/Lw+xDxNluY8zRiYGbfjWOwxbx5klXwwDtVO0pd74m2cHoN7xtHhBVT5lmk4KajGz59fgSwKRF
9pyLJBcdYLGqYrS09Ul9j78J7CoSa/gxdz/ccBLCCtbxUoOvUapCFJkVpbsJM5A5zTWZhmJWWV+d
//ITvNFhhtEgGRSmy+lL77IGmWNC1ahcDBro6n5AJUp3V5M/NgyRxypZkwhrGasZSYE8fISszk8F
Es8W7rfotrdSb1SSDUbwKmTbVC8iFQ2ZOjdzrfyjMTGetymwwiacH8z7kyIy9GhQj54jUAAZ/CuB
HHOlskYzO3vE7pAY1mSOZUCp9CT7lmVADlxtHyE/fU8O827nqcJvz8u+GsODAWuqqm5x5QfA19tE
MFXlUtVg3FULCeBnbPHqDDWS93asOVjw2weimTKvrBLcyMpapAbAZtYy5T8S2CMLUhguKUTLDlZA
h3R+4NCbqOqqXz051nOmqQIGsjXMqhDp8CJI8M4be0YV9H//Z6itKguXFYkaZNa5y5bY/08xRqF9
f7Zb3s2dpEwmuPdPvl2GndyQbTs6dfgBwCWIkVMZPhYN5UUKLLY6e0AD67xc2TTHpaqYS+pnHay0
DNSEcRWrU0Sv3+DwlR+Whqz50JdSyxqI87SuSOVVZCg3l+inM6VTfzzfMfw/aGWwUQWV1m9LsjtI
mvq8lMcZkJR15mWe6arR3fH2Z9nPyg5UABK0hPNtkRFL8NW8LJONTxVgIzu63jp5ZyTMnJApZPwb
dW0Xj4FVI4H+L5ycSsVhS2fh6guT1B41ukM0EHpxBZP/yeTeWKlx9ZB4k3Hh+Sz3qLw7wLil5enk
FUfxHNqCUmTTDXy5+HWLvOSuE4xoqqaZwm+0VYn/xMVju8q3F3TIt4GQXgXQgCssiEdxZcWsEKLc
xW4HT5VFnck5qAN9yfSEgCcxWQCq61Abw/BZ2+a9aMhLxep48OGGTXcCuFUeCZBTxb8FzBGEhR+z
J85MfzbMv1Ruz3Ronf2hN75+9uDF42kJ0AAOc0fHYc2BOVsQ8OCsClv1bEKpk1iRuGHchTlbvvOX
683cfhGsRVs0LmCGfnG9xiY2Fky8HkXE8xvHImf5QTvOIoBPTHGFgRegaCQ+XkSgkbyslVFcx+WZ
dcj8XLBN2FXerv9+vIwDPZHK+XVSIArPzSNVYkk8b9jvmNS2w3DWaes2O7qEklUeOwLIlVJ2otQ4
ywP5NgdG38nxCwoHaODimU3eWDPIV3eodBWShZlR+vUl9yQmhmhv8O7INfU9Ucnlec/0fBJ4WIFd
dBXlrddtL9doeqYih5ZuhuYTaDjQ72djzd4YqzSQMS14WrV07R+FNttWIbc20dDanomWmDAmE6tM
pLPirPXmYRSXtM5Kdj7+t4trbblRwLhFRMXVri0k/oSzKxetnxdjkuNWKpgULZ736os650SMZ6Bn
nFbDZYdwcKh2a7OpruP63ZfAwFrzgzy9dXUKjIJcjuvQu2S80IIqDxxhMZgb5K+O9aJXdG5N3jFX
YWnCAFBpghxPYOvCRp9vKt12PZKJZc5dBOkxK/LIR+kSCl8VtD3NFnVeRsCzafu0/BBtnZUui9U4
YNDh/8Ao+QG7qndQsHaSU1tJcl7h45wkLRXdrz2XiC9TlAJUHtq1dMm83IfCMftNMyEg2VKAbg3C
dyGyEgOP9gUsj8ejEaB4tfLdzll9zJjgAaKtWAkJdqMhKJLbUBqFTl7fi7qOQKxfhsXyjub0stf1
HTRvucg/1e/aSu3llfqENdYiDJQpA2hX6pMi/hfEro7/4d8npQPSGsTTiAE0RgWLCTxCA1d+UW9t
DVoFwCjeSsZmWfamQAH7bYuIGfXYk1YpQldX67ovqvb0VyPMh7hoi14cXbRTuecE7sXJeJW7uR3v
2e5/DPVC6P3ektjoHmTzB53ll1iXezBefjHUtxCmrZ9OC5PwB9gn2jgv7czgSlqrQ/AMVEiZnUxl
L5OAeYC+60XFyFOvcPkKPUL9vUGb6qZ55eApZoN7/sh6+liV/dZf2MNas4HC/7n0MP4aQ/Hu0HSy
FUSlYfXFeHmQk9d6frEgQLdXJaUVtLKpOEBwhZzau1j9sIfg358fr2bTgza3fvD+PeAbmkbE+LHk
m0DGGPaDP0Tcqk0PuQ/s9yW6jYK0+WH32bXmKE+NfCj0luFgq0YT9dH+GQU1QeGs14NVxBnu6bBE
abcyjsjKnyk+FWlBMoS+N4Q8aF3PhZaAs5EYBoYwvAfqm1lFIBPSYy6EorHW+MWOeU3aEEwu3rpv
HFuZaICp6COWj8enRYNZppDkoZp3VLegY38bRtGLJ3qTYQzPQQHllGBzObWR+0d3jyoZ/G+XYZZ2
1JLFWUL9t/gske56s8KUMAghRCV9HXtUrg+672hT3kom/F1hED7QmnGgcY8LLgzWYRHk1ajH2ptE
pcD5qh1WsoDLW+vHUhNTTtRfd8w+WAGUjHrQz+K8dJmg5U8gV1GP2Y7ciEuOQhQ8bjjdJWSNMX65
8VAiysbhgq13kzYCekewo0iYq0HxQcvTgmahtyM5KBRGOwtTSgxnfuR+rPparczJBMNjFrxfNNkJ
6vrKMtRKudpS2it2hiy070XTTgt8Dmq0MXka2V2oqpd4IvjtJ5iiUZLlBnSWEx1zUrZQ1cm4DBS4
Qb3YIzXX9AoE4ga5YKYdxk9bmp/UPSK2yTa1VVI9Vrfi0IwhMqpQDHIbKDJO8bLII7BJpPY+Fa16
BLkwsUNf48q/IDb4PyLJqHoLHRUASfSKbnlcf2bE0VLdjlHxA4itAxncvz52oFuEgUofZgjGXXDq
HaRhYBo0u3MC8hpuOoDaDj+fD+954w87GxFdOs6YmZ1+VqjS0zpSOxYnYhQYJN/hstdzsL47SDea
SP1r+IQRnuqEExa6mD74LGi1Z/H2WYUib7TOQVx1a+/OBzPZY9OdhpaKHZy1zEEHQtmEkJ/xCrRx
LclVDxO5aFv/V+2MvJWK1lIOSY4nocu+Ruq5I+t6TWL+9VvJDtrj7IFUqe8pPvFgGRMCic7NvPYL
gLN1GINWTMV0Qt2Tg/NJkDLR4sqpqSKw7OId3Qb/XFHAh6k2u3LCjbE2jPwBj0q8qXwrDQsUKOiE
GVIwEGDvzf9SxZHjXHyiMCKXiSNMAXAvBpyovxAg7lhhSuY0WfqEbQnXoiyR/xInOAYX4FuOTI9G
DEL1KT4N7mFQM4ktSUI2EOS+5zJd1LSLmNOm+1cqQL1qk8++9q+MhLiTqoB64NmrG9x7PFbXivZ7
J4tlyHBYPTGvPB1YVCSb+4yzy2RycjnvykAfXSGxZjsVU5S/KViDwINIKYRW+TYyx8odqYrJYtlJ
Jg/yqam7P+q5P4Hp07FpWVFC0iX4ObmpXAlV0DbH8RyK4ruO3eod7UqeV/CzEaC8rcayda7H/mWo
gvuSgaEQL/ln24BXBgTb6fPWvxxmI/gCwC8+KxHTOAh1NFld3iOuPhnPvFo8IajjqzGDoFw5xHqB
c7nPB13rf7G/X0H/NXd13TGfmSEp3MQVeGQCwhQPSDx7QYDAbixYFiORtEBcZdW5KJz7+6LLljQw
kxUFOYaYDmjg305zEJAxoaUw1sP4zZFmJvGOVrX7MLN/JZjnNF+BDeh/YthM6Y9mwUetP/j4cjjP
6Nv1sFQNxiFX8n/bjsfB8mabbp1QcdcaF6dosSIkVHQhNqSJcAGu5gyFWTdxeDXXDp/qhvMDMHxf
NQEA2uBxaZz8xTGCqP9oTl3lJGECcVoWskfVdD7bRPAN+bQDTsJPtHq1RZOcQaMXsqXVuffig4xe
tAAEkXXzTWkBFAT4fwFjNPDt/+u6WT8Vk8H5J7DPRgumMmq2N/0bwBC1h30dd1wVIDnOtci9h8de
mKTk5luWZqzP5KuQinqEp2lG2/39c2lyTn4OEf6bUmJSg6188PquIu8X5zl0EKkd3cn2De817wG2
7bq9NWbYYKzpQlwzP5cNpsLWLtkuZ0GEuSsdqP+tyi47Kmvvh0qV3OdvnkHYTCKKyIeTjG/W2h79
3JhbEgIENDaL27GSbXGierNhOM7hu9V5lis35V8xpJuRnIocALXnE240vA553xeWaH3+64h7/ozt
UNpeoCU3pbYekD4MCsp9gRtIEUFL4LayDmy0h2/wOak000IMuhinTQgStaHjPzD0gTnq6y6NsrDt
onDY7JDOJWqqqjtqE5soTwZj59BmFMmqhuWNw1HCmtoBxnivOkdZ5hpQhjiknYVXPnQwRoiiM6lI
J2pwXLLP38plIItYkP03ruBK7JMuzEShn5xDCvoEzQR7DnT8X4tToHOXXg1QtRs+FMlhvATWH+mf
d/HLXTMKyoN18IzR/gnkoL+CkT2WoBWAPQ1zGjqH4lbzUTszlnxhx/oNAlwqEil0Ojybs2VyCtNg
SohVNhS3vMwOZgUB2dhsPUBBcIFKgcBEN6aq+3NiZB8IEW3soTJLBKSuwechoU6RjqLeYWCZPLll
F7Cpy2vf2AcoeqKX+SDt0ERHmgFMfXI2FkeDrmXNp4dqHT31Qij3DlJz4URrIi48o/MnsLTbay4s
f6Dk8uLSPGV8bl/qdysY1n4Tcwf4r0FFWrJrMG8hiWB2CL7cdJzqu/JDeNYlK4QqfWoCIf3eE7Y0
mPy1znp8FiQL03mXw8AswqI09U+naAC9rtqMaKzKoEn6R3DrKqpREqpzF1pncl+bkX2idXCF8YJT
tI+TgorZjnIzhXKMMp5pUPXq7aCH4hk25B5kPjk5rsfVQPr5NEE7OOtvSzfJQQPKpFO8HM7Ak9Tv
VRpldbnvMbo2mBgfKOQNX3fefC7sJkVEhbt97ffo2ps7kdYXarMB4sp1jAPLFnovbwwx1nf+I6m3
dXVOtsjUwcB5tmpctXMbzeAGwf8AY3ecisH9DCHqQ0sPnqhs/1ZaL/OjbTQl72zCOzIkOdy+71uO
GP2YOziI9jd49J++qqOAqQ+jARAXzKh0Se/Mcd58TF3e1EHKsiNj1gaxcUNB7PGAMLT1UGsVSr/z
y1N3WSpcuUiC2CvAHBI//y7sEM4hQxQJiJdAEItviBpZJM37sUDAAyJVU+k2UoDmzhIDF0VfgdNt
XEpKjC0Dn5uqn8txOcrArTxRSDrqEnuK9wLwB54c4VjrI7hKLTHx4PhCHSvYOqNadgtOiKr0nWGi
EK5iCxfEtLfKasTHNqdHNjYedYHezAwjMuXNOylnuo5RcxNXBsw3UX1AamYvNN7O9MwvTD11YLO5
izWtIb0pswvc+HD+4zfYqhRWw6CfCrs7WNUE1GaLggVlDfiLoHG8KW0fTb3v6KKLbuuCmSWENR4k
7Cu2LHBPEELoBVRZDvlajmv/pIXUMtxF6bX0WHUOxxlkz0cbhgWf1J3JqgeQMz46Sj2DdMt2CmM8
y7G4fuD0KT+dysj6ths24Ue1hmjbCSlikTJeqPKYHgZ3AiLjw03bkjZvSBElhbbqmEuhcbOY31Ms
h14yEJDxDPVK5TvgIbeNCSKEAduQATb36gMCbe6lYowX9atUs29QUMU8ezwFzBAumUQVDSc8d3HY
N56NPuIXsGrJhg67HmL1Zle4er6177tC+V8WNRzVFcn4UTAHgTf6wrhKO+fcAiDBH5gx4u0yS5mu
v0TwIBseLXItfyHdllWTkfWlxdC06UvRyPRJQCbBeboZn8418WLi7d0COxXQzLNuGqJxqqPa/Ss6
zgEyAEzbpruevuLao2Xt2LSHzM9X7SFC2qo2q/cyAi/lj8uT7k+uKqJzjzGJEyosFrDQb1PUeBL1
/aHFmky7sFvB/Xk3uVz23tB5agsuYpfBJHTEXhxluSvRY90rw6Kz6dmcTft+df7D6Ndb8j3l1tpQ
r0JGGzliBB5CWw3WUgp/2otEYkq8j6Z92GYyYLTMPmOOEq3igueRDHZueNlcf59JTfs2JmDhqSA/
0QmngMEdgvm+qYhRwusM0K/TokS7M0vUccOJNX9BsuDajcoXZILmf/+svSIUWwzgg0ojk66uz3iD
0kh0yjfEuPQJI6cpnnANpCW8mfZUXK5BkmeqxToF0QbqPCEtGAWo78IMvLk3joLdwJABsLB3dE9O
bz1s6RJO+yp5aec42VIlD2ARnX2yjcPaB+kEjYC9rY3v/mW3okSoZRSFju8rklzCgyahczEn+m3O
eFspUVOPrC2JjPpOKK977n82PlT6nXcIQDOVdXN2553bFbu0U2PFXCjC9xvHcEt6pIk4XH5yxv40
t2J4Lnf6dzbCzlG5TXeFAeo4jIUJNiAZu1u8l8le4SladKFCPmEo5vDT7AbvZnLTUc3FAeeB2O2N
7Eu1Q05w1xBejCUjgFgbZgCn4p6J+IvrDaGdzynAVvJUBT0WY6sarf9hOWHjwsOYXhG2SxD2tTa7
vm9wibbhEfJ+BjVtWkgWSDEtDMaXUpo/4PLi6P27rhMcRp6i7XOo3bv5Tgpbs9f7MqG0yYeTiUjF
Tj6MROGl0AKQOe/YNvPvMKSNOQOo9wjboAiq4sHgiQrAdiITSuKPRpCif7r96zw1tdCcm05UEDvY
ClOu1MeQiX90wBACqzcCkaGSK0ubq2QWRLcFG4QXueUlNrImQ/EpV65HCPftytYj//OMslRJXvxU
rMkjOlERtkV0EbhCHcYk6SzRSDLO6BbVhtYC7WfNbPHLbiFbGFWddtB+Za3qW2jAIN4WNu/gDvc/
ZCiAxuPGE3Ztd1hfPSrp+Oyp1B67R0uTcRxNcMKpMOOOI0ATvU7wg02r3CnOmgh3IhJetqaRNUpN
2rfVPIfn0iqPlIkocGUXJoK6qXJOLyLEY1BevH+zYwuIZ04CqePVVf8uI2sUWcxC+6hHjacM0HHm
zcOUld8WMQzElK2J/q6OkRz8mWA28cag+c9ANttTGRlEJmYwKcaMog8juVP4K+CJOfXkCYM3Djft
ihQurk70SrP3OktE2hfUOKtvP3bJmK0LdzFY5X/YA91bLV5dcCg8tVNAwabwMjTjGANDJ96XXtPk
EfaDSt/0tZu6w2alRDyg14SH/8RBV11/4vlaG+MC4TteQq0L9WJbFQbMHKie6AgkGm9+trnolexv
ipOPKXGmaosXovG3rdqZxvX/yj2tjMAYYPIbuC3PKEBtRpAUIHzfIa+t5sn2UsEtVuIZWXCi3OqR
A/OMHvZ9cuvCoHOrIKAFBSfiKr5cHzVq1/inqr8yM7WsZ738N4pulSqEEcMiuXdQ4/GWMoCbFFOL
e3opT1mFfSlLv8724S/Zm2fyDHfRN5QAf4IfqHXMeUYz4OMf8+MTdOrn95bFzV57gTGfSm0LLXAk
GpAjEGumk8qhGhPLrXuG66O17jRROtaLoLaOhx5XkIk1m4F8GZiyGRESb7mnt7c2yoOIdLKtqR9q
sO5Xj/4jl9bPhknf4V4XQUOpzYW3o/FXXxy/FKbsBeOa1ztOaV6/wWYQADS7pRnBf7QIaEXlHSey
fF50OIr6jq5Ezr3ZZGEI/BomwVInwcHoUmohIy/sVyVt/PZBeHcHMBiWuKLN3z35p5ZvH8mlnCZA
COIi0ZSDYxJ2XASW67Kl7Zoek27i17d+7Evsto5Qr9A6lpZY7qPRSvJ+J/Tfy1dZwaKdFjMUe7OV
0lRWNJayjTAFR/kyJt14SVgW0zK6VgVfy8qrFYHzQ0r7LGTBV2b5ND98Z05fd0mmANMiptsYCYaw
NR8h9nzPqTBK9Juj4nhoVA0JzXpCLz8f9k6S0yIc8w1YWgaVeTn4iY54dyv5oevWLjHTlxzHA9pw
jpr1pupXjAw4oT919tT+4eho64Sc+X8u+V2sX04VXp8qI9x+T45QcOYJMzdjmP3BKeRTUxNWFi0m
EY6qxaAvzymGoZlytRVns9OXcvr+dk1CIYLKQB2qMJGZXWXwM8bcF+mrYl6rUHqunz+8cXi5Vqok
DFxSeWMSs+OUcOZ+x8Xldz4QYJ/NSXBuvkW0okhOvXiSJfVUzoFQVIIjVFgpe6baZD1Fi3p42wgM
wnxRlyZhFOGp1VpLjM/MFoblmJnRbTNz6ZMyXwlO4iLgW+F9GPXCZqQeNsxVqIzJkvkCRJIJOdcg
9Yjp4U6URBmiGYALzNakW6wND+4nqCzWmj265AjhoVi2C3x6aVwDKGuhxDIEAXeP9LuXjIilL3Pp
7SMYJfwFPXThf4NxA3XUxuICW7IiH1bIesYO1k8F6FMtvdwnvGu5ebD2mA43wqCZYxJ32iwgdFG5
ALyAru28ynOqfM6GZhjFbmgeM3gcHywBc59MfAamanzSZd4XLgT7waEyc2jxZB9oICtNYprZbuJs
BVgyu6Dz4Cpei5EJXFbruxz13cxCF5MPT2P6+zcf2KFp1ErNa8fyEm4+05gw4FJs59M2QlZWEiyF
kP6TpnUo2/bQKSWIqi8TsYgOXLonJrRko3/oFjsNLkeEPVSMYU6kY9eQPu8GvifYhsgYAsV+mFL7
Zmuh0gXWLT4MkPuUK6i3ogIMTOaE44sM/S36BiJsMh/zujLDlvvuifiTtRVRM6Ejy61tXAXrDOMr
0zkQOkMIsynG4BgEvAsVAv377jGCelYqhm+Lfwfi4seCoV6SzqUBrjr9snCZbXS8I034hhHlV/FZ
SWi9j3RbpOs1tykoRHWU5xyXknZ27VP1Mg4K+Co0xq6RF8Ulh49NciM2AbSZFtRJO4gJ80KR6XkX
Dwi17skiMAaT7HEUgO2S9vSOn8/uWz3B0NLupApIJmJgnYfrZFXIOR3TEP65ARJ0w9SXVhvMU7RO
DtIm4xmDyaOSU/Vnbx/7aWUzUlQKEQcwAE3reJv0qrLd1e20z39Q84rm3+5f0+bNqCLWZCj6DQL6
7wpAQWezxh0+xOBWVVyhkeLfuvK8WbFw6KAq2jChsV1d0GvG9253eVqhC/yQ8wuMl3OkvI59LMhK
GOhX0XDHX1Z9JB0cG8NSn3xWDt8PPn96/7sS8HmK5BIwxbqP5/2iVHX9lXrsm1Os0HffQV6LvL/5
6rprLiUeFaZ8rmwarflEj/5itCfA0tn7nzr7BXUnM9TeREa+5awWlBykMIBCD5mE+RbVPkHDdt9v
2ttyvfSAtizvNDfFtQbIsCK+wdpPYeiEMbzB+Lj/4Sbbcn5dRb89wu+owR68jBOChugAkn+laXL6
13Gh+0nb0Qgjm38tSCCesyl745QNm+29vjFH0ZESoVdEMo+nb4/APwbqKWo4qvSr7dKT0D9XJs2d
jLAiSprlMfJQjQBk8t4KpGdmnKMV1UwPdaEr6qpFv8oI6bEhEkr1MTpmprmoiAijohjzHi1m7BlT
qjZUlNmPmGyw1uF/4WzxbET8EefRBPh2qD4a7ojaxkNFkXx56A8QqkiaPZmmNH+7Yks43BsQW63A
VeUcDtjQzTQfLqiQgoJK6kY9/Pah0XWeGHh85JeGL7IzNbZI8Q9dzx1Y/C6cubh9g0QVvtaOkQf2
pif9gW0G+oPqveVdzsYUEa2t2VtfyqHu+zEs8pHGSXMboexz1YgjiNCMDCiAsRmfwScbvVas2n3Y
9Q60B77Jk399w8VtH8MGZVxxaRvnx/I1NAyLfylb2SMI++YqPR+i0101NVP3d5hi35Fu4B4g3sWf
C7uR2vNccS+M0s+ldBoPk0O6uvcB/yDNQFv1hZ3ULg+CjMfaGkcy6Hswlmgfqew9mpdKf0pYlakF
idUOoOD+Czqwl/C28OuzWGu5JV5fCkL386pWqTYAB4e6XQlf8gUa2SB3LDYwyVBasLv5gwMn17f4
KlTDYz82bf+skmB+OJaEV5NxUfvwMgXmQ7WThwkeVxeoVC4pGD8dhsOWx30bwdipZh3fJCEJ5HsJ
hmGZ9+F4UJjSjwmp+CGQKSmFGpeEkGgj4aXomB/j0CtHS7LAGRUT4VigmlXEtjQFvfQZ982D2uPP
o4HQMO63/DeA9jkI1Ua5KEa0JLO41teB9/Aa9WcvCzZWjIq0IjtlfmgbREMKN/DF3wvlLsmgd4kn
0Ic2nc+G2JIKq1DLd7SoIWCGlw+pErLa0MRT/vQbv/z5OLLh36SyZGh/vxQPy9yNFiUO8iTLjwdp
UrSiADBGxdI0F2Eo7+m2x7BJis3MGOeBttCrGLem1wUhUI7wrLGY+A/8WKlncuq1Ay56wUUEFw4s
IMOQZXdKQHKoqUUU4XjIoSFVCEIt5WE5Wkr9vX07Wa8Kx5T2WIYQ9xfTm865Gi0w3VLVqRw7Dsqz
+6aalbHNKMbXzN2WV4tCy77LEKU9hXDeb5QRxlbXzweLW/t+F+NFtubcMQ5EG0XkifnEOWuQJ771
R3HmbGCqihP0pMA1hIRhGN+ETHuKcAYmfso9r1gIhUf7ZDF32DWapvTcc1H2YnFzM7jrwUegD4iE
y0QSgaRlofmC+yXnt46K0J5xGlmZgpRpYEKqqQYophgtuoNChFxToNJnYSHOYhHBJ2jUzySuH3hK
ur5f8kiqk1PgUDhFAhQ2L+cK+BK98PRN0djqVR8h74qE/AzKr94+NbuOoA/a4EmBwQbqn6XDUfy5
704mKsN0T95DFqBBNvdIvKxY00Tw5rEiuQgljq2p3kHsMb0gTruMv0D7w6tRcIJ5d23LgYia9bI1
Rs8UJ2GReFEnCpd4n+rS/QRHSqWdSf+ulcUfFzwUDkvwBs4A88hRhyYfzgSJ+jZUeU2SHWjU71c6
VHiCCSzxjoQ8POBDF67Dxiv2sVfrolQZ6T7V2AEeW9ykjnzH4d61yIu1zlVndJkuLQqAUMP+8qBt
eJ5QaG//ocx/t8L3EWHccfu+7hi1aqXw/Vawfd6gruUO7S0/NL9w6Wienz6XE8aadMwmOFG4umG8
QTwY3thWlnfrODZTOcvgYKgcfo3hAf2g8bqeg9Ex2ylSvtCry9hmWvSzQPhrpjdbVD4zsSM/5RXv
TQtDN3JjOOeUaQjB269Nv8iJ1iaeR/L3HrQUKYkTxWlFHuEunV9HU4PqCeMCoN+WpXj8fmGxQ3rl
K4yhiIsd6CiQrkphun+ug5kKXnymBb/otOxz3hOkJl9qZeG34+P1CLVsVzH6wd0ypBbexfRSOj12
POidQ84PZqgqwv/1Kf3jtQZEb4Wuy4IOUIb34tzEHRjRbsgSloPH5wvxeYYeiwyM3ARub3QJp5A4
oiqsSUlvap44hm1w281K+EQxQ/MnaQInI9tj01XNZ2uAdA6jcaAisDLpFoetm6jd0x11QdZ+HOr1
buA8JW++ezoihS5PNO/FvTl1qn83XKDUTxtkBI8Zrv/kcKc5VUjmgDijNv445WyGSD5GlsZcciL+
3B04fARhRtk3PZRbas2TJM+mkrASjh2t1pYJdjXTkcTeWR4eNzA33B9Aa3ImGNHtVUz68Q4KvwWi
tTvNF6jjPkiw/1PpfApgVWnVwtSR+Bth50rRhABekoELm2Z1V32io7khQugQ4/3OYw0jRKkoMItq
Fz4sD91//TQNGYJi3MlIapw8q/GtxxmGCiiscYYy0U04XL+8B3yMTpgtku1vs1/H5FafU5r/XWM6
P44Cv3BmhVSbXTEQUQwJpdoezb4gR0OlY8qrn5uWz05YfxO429HqL8CsMVm4JmKEOmV7viLpYVVW
d1GMFZj+y99lx+W4PpCas6KzSkYycl+ExwLebnHre1399QwOrd2iEbM6MiPrH00fzZSq9ANxZvjo
QD4QwQ3w0qkaqmPpx/iS5qOPcE/XaLEkjRAE68zGRv94Hsz5Y+dXFq+sJ8iamZjxI3tNcAX5IYsr
hlyqP0JBOGd2e4CG8cRhQX83o1dKoVPbPTugE06pKCZrvsdnvFC2Vbps156tNc56w4SGPWV22vAO
xyz3Mlw8xIyqCPk9X1mu3QLivqGDGIrVAlFv3i1no9idhGhWq+EtDxOJEJMDOv+sqq88F6r6awCr
gOWZkqvE+sNaKyA5vnlTM3nZUVARXWuT30YgmOffdHyNfVlZJrB2YRngpqZi+NiOov1lUZ1tYhYU
ZmuMYTJ4aTbVewRqZ+DCee+ankaL08uIFtaIzyxhQ4B6c+sisBaIPgMGmCOPzSsYHJWw04g7VIlU
sH/8zVIvx5GBVjYLLhIwlzBkYNnUwvcd48mjtB7ZGyEo6fIELdBNCvzJhCfoflFLovZO1T9y1gOt
iUcgXzucfD/aouxmJak8pWC/OTlHSqPgVS8gcgW4vXLE25PPZIZ7CfTakLpLU6aGjEKqVh/3X3hl
sGlniPuFOYqto0FCRzOQMR+8LdowZZFeoQ3wGiq0imDrYUNCUSYhhh0poOH8L8HExvHefhJOzQjA
NVS5OgG6r7YCID7zRKsjrSuVOOBuTw5tLm6/eRF7MykCdsPR7eKs6BvdDZy4XCLZPZh4YkWUKNbz
ZenQh9N77Vd5sJAqyMXsXt5caJjUCp+TcI0DXQT89e7EG1NnPOW6K27vkSSzSkn1C+9KHPg31WNz
YqzG0YP/JCTFfQFEJ/B7almYrMszM7iCOR9Wg5Wjz4aZDevCffznLYz7YYBx8Uie7vl0iphpywL7
7hW3GDKzx51jQzR//orI5UOryvQaTsvOKnxUsrsDHlntf8wHoyU2y72NGLYA2OszLlyH1zEhNcUQ
5yDQn+4oJY5cy8P0jOMFIFh8MOzPsEKzaPy9yUF49s6r9EZzW7dHE36i/vaEvNqFNJmtHhAQ+uT/
r97D14W/fSdcdAB4a8K0CezitjHKtJbL39EJ+1BOnvsQBX4O84lazYrB9Vxw1PfgUVkuN8fQmOnF
Gg63SCY+2qcaeh5s/6mrokF6LQ8J87DCc3bmsPQvL3zIgD4S/FhItjhEP0sQuWYkK4zTrA21Wtda
UyeNkj/cX4M4on9KwB1lOO18pQOs5Y8fkqtDcvwZBKR8P0YKmxypBdzY+wlopT9eBfB99DTQDluR
84oQ0duv/E5Qn+H1lYEQIzyl22HAQqVMByoJxCDvc3AKZT4LYAip7mytMASd6g73b7VnreKKiAbM
6dilCyoSlA+shDVVQgsBHS+k3QPiZsTD6z2H+2nZO5s87zvKBiA/MsGdsMRZ6oI7LysSguCiq/Uo
6RyYAwAEEgR2oE+obvZ6GWjWWQV59W6dbUsrteWEU+q5FQgRUdgULDTh3TbZJruzRZaxcSUY1Pyw
+gwrAqXgpcV67mSvL24WdkPg+HykdpxzYmvpRHOvXJ/dYs3GLo7Pdi+DaaM3XFMmOCmiPA4ijtZ5
WkAQr8TYrvVHblDCGD3Ahn9IKYodqrOcXVb8nfEvzIiQNKy6zClfSv/MhSKeB7wnTklmL3qW/UAa
u0yoBEwJzIjYjJdYQZvvhCLGXOoK05beZk/3fscoPiilOnADgkFRY8ze4C/6KxJ/+UiCF1mwH3Pi
eBweVDElUqgvxBMO/LEYbU3cEqnwqCyhEE9mP1PI+LN3R+XRIQFkxbgA6zh4I7CpDfhMRIt+JgVR
zBZFFqU9auhtBFvLyrvfpXxcYjFnDDC8eSgZjRYlIU9eOtRUPPab54hH0e/ZMNsLGFzWxWtW9fKF
CvbYOcugnzF6KTM9Wc2Cot6ZHeIDqD4MxmsveDubcPAUDGm/1zU7lw/XoGXybDJ6K9K7cNdIHEs/
FnAMa+DLF+1Gab730s7XDRcTV++GPbkbgMPEw+1lXcUtDcISZRLdDzT71w62ZAcyjNP74gpayxlL
DKs57JrcyfRbu3/SRhwLYu9bNqZCohYmPeml3efBglhtmgfZkSYDJnLulhVZYlisUx9c7cSMOeZr
FLcoKzcq6KAbvAcD49hV79rK7fVkYxVI2j8IDEeY7aNB4JFx4iSbvalg5DP49o6+qbAi2Nu38yoT
kOKjYzvoz5gR0UOZAFD/RDRbMMAayj8OfQbqJj8fVqd/cUQbVfKjCKA6ww7j+EqudWeVHkSmIuYY
k5IZjxJf74FqY69uoWTdiNkTArW7VoqSdhgFYJV9/+zi7Z1R4whvx/Rl1UGa+EDETei0A9ceSWjb
I78NzcmFPZLw0t0zDVfOidSgzJAoRGT2/EkvaqCP8Lk5qjGciZmq6kzgCRYXtndQNRe13cTnG1+A
oruxTzrWtaZc6+mPumd2yUpKqXZLb2WGgxh/keHtKsd4GY3ltpEBbScKXKYm7oKeG0e45YEeJaw+
y0tRtFoJLHVj/sptChqonDVJpm/oy05Qhvsl2Dc79U9Cw/HcE0oi8bfWHsOKhwzHvXnTMhFSqzxc
ZWwcWKJNwNjTo1rfrqF1llDktSAbKK94AjevUnn1itm9iodZ/kf7zAz57uKySMWwhKpD0LziS2Ze
0e/PP3xTyEOhXrWg4DUKIk1WkoFq6hx+T/wXNBOhD+4bd1bby+vk/XdQuVBfHzx/HTpg1H+P04MV
Hrly0RZUCxWlTtJCl3hh+M7D6YALr79QQmYsAuwfMZ5MFAOQ/nS+dHIbld+Cr+BTJ3rT2tEka/JK
sQkHpgpefX+SvFs5clQyyjxatYqfQib+eCGt/vQpM/fBO8kD38sg3lL4T49mZtLNqSAsxhun6xnU
SqfoE0N/yfrcQrBeWpT+fYpJj6oEkbB0k0lxYszRIY88iRUN/N87OZZjCn+JreYokB9IJTpLnY48
+teDVWel1sdw8hGYQnaC8VXIkVu4tiFMhEbUl11zgoYwdutVf1TBblYxKrj6rO37BJYi8BZENQJh
F/Y5wOAN6R3+Klj0pImrovJdMkBSV1kkTMif88IDifkr/pcQFShsLQdKlOjwEgxsGgBfZ+y/zAEI
Er2Itl4J0/jyV4kqmLPDAyVXQKy01UeFP5geu4vSwMfn+AH6z2KcZoTAZeadp5W7MVRvKJUPDMxl
hCGtp2HD90fmKGSw6jr2ILYNoa076LmB1OpjR5nCqBZijQSJyniP+xT8hSgtjmwIZ7iGUkVNOqRk
QssPnwAvLadtjC3j2S580gBRbbADJ2BhaxBam1UhYrIkj1trLnTHIt33dB8viomLU5lRzJtJEV2q
s09TrBXPi6IgVHAvAr+hqbc+OAKBKE/eeYeGyRxt1EoiwyOPwSl+shgNfShMYuMyB9yvUc/rFt5k
Z3nJgh4fOBnV8lri05dEo2Amqdg9T+4Vxf4cB/sAjoQZCQWJW/k69p5KJCEu9I7lFMxKzBP3DG3a
M/rpAsoun9RvVo6Y63fZpfmWNpY6n66WyWIlN2rRvVt2sPK7fq7YapOZijgPoQxOP2ZzCB43n889
0x0BqTB1TW2+fEANroirQACrCpMY/New7ABVnfG2b+pG9i6tIdNSSTOWFKMPyj/ciF2WzWK6EFJJ
ro3EOAjm4wxdinx408U6gK8HK9Ud2Hrm1cshWORcSukmHsn9fO9FwZp1OvQonNaHEg/hU+PiLqxc
ZFr+k8P8JxN1QKJtOT6IznSyOrXBTIGBQfh9Aa1fjVNNHIMuUrIEsHtpkSADxkQML08b6+VISSFZ
SPFgBGL+0qPTlr+17sFU6tb/C7mBl8prVyJ9PA8Bsl5Hb6P6OMXasM0K506Nb5/uRc4pCmBnaoup
Q6PhGH8NncG1yhxJIsTrOQD9wfDcjeNksbEZNN/Tvp0A+j46OrXjBAP0Whkbbx+MUHVP3xFicozH
QRwPD60GQFBn+3s2D4n/PM/Bvs3BZQuyAhr/ei3OD+7HwjGOIthO0RwrTzE3WC9nmG378pNnGVBU
Hjn9Qr/IrN9/taijHRYbjrOeZp+Z1N380SQe6oXdTq+CYecXqImJUOxM5nqQ3L2zqwRu6z2zk40h
o0LaVOgCiDY4VEQIx5mUYWFxAR69KsJ41Xnjm7PVK1gFJB0f5LYz0f2+xzqp/JT3lILajI96JgZl
mRUtITgIgCxXc9Z/SGGETg2R1vbFepxgpzQQtuoCn2z97V6fRlMF6T4JuydDqE1AcY1uJ9berFcB
8MpYW8kQ2rIvwx430wAIV1eHfY6h6ftblglv3CVsUSAS3wrQF6aTJg36l3y9m5zzUIurB9Bfc8Y6
f0jcHyfXl99ScAH7b6QG3KpJTXDtrSFBvwDDeGkbDsqlZFVd8jwYMqapUVtRtLeo8Cz86qaNMi6G
aEsfW5crnt0sHadLmXj3Nm/zK9GdzcgiaJ7H952Lmjbcj7U3rhFDmKR7i5J0Cz9hM47VD3fC+9PI
icPJ7uQt/jDv3Am+Y/UVUcGcqQ5afJ214qmawDVHoqcLjqhW8fE0UHAZeQZFwKKmqb3mSavSVOV7
g2qmTikZg43KjYX9Bke8pNZPrQwdLmOzywcX4mmXpEpYC7Z7wYc6Wl3n4sN7SHyGP/6pE+bp4DzH
65H+QH1hQpV9iZUTNQxPu4e7435kmWWwpSBD+Vc1DhiZleZ1T7GB7vhVnX0eyMLCDCkUYUznAshI
FJnUd+G8K3tMyVt+4e527Cj+HcvXiv06/vetwBe3V5dEiDQ9+NRNGH3vuqvxY2P0+zSD2O5o/OXy
gPXKwhA2vmL3v9IQzZ9U6xHfC1fyzPRl3Efgtt9UPpMVk9uYOhwKFvEcWGKEvcafTJjhbeyr0xhK
9jpzgravJTz7/nhEHdtyEdZS+bo9ReG2Jf7kF4VRLpBfc643ZkaZSGmpzB2ETUneSjRfp+sUxZhP
dPLQzWuZeiVlSuhBzMmmps3rw2A3rYccUjMpIV/B83rYd43ctDUTfAtG7ImDOlx9lAxX/cSr5eD/
luJB+pihPwrWodYJmK88GlqiQaH5PGUvx0pvxVb8TghzlT/x96gUbJdWn+EQAzg96nBQHMPzOVB1
B6c1NtNxTo4Ad4b2AeEK1IBBUsIiTWWXA619a8367/bSV+vGuFrHWs/OMViBQNSAftA/zhvvLEOc
yLcw4iatudOyULlo87ghmgsdmBvIaw0IxLJGwN49bboxjLFKa89d+LSjH3QoRsa+eoErGS36U25M
LKHXPiARoyDTttUeIZMEnuhWFc4tmXrpz81xuVfqrYoHmTOrDPJyVTNfHXKKCEIoXU8q4MBshONB
6sYxlDs3yJca3rm71/XrZj4YQ1q3JtMEC8/ERpAcIi1XTFfMoxmS+4NW4vE34PMvnyVReg4Q/zCM
z3EgHMG+J8VSUT3upPi+PxMFa1jwW1MtCI2SC/EIj9CZqOnC7O/gsPC2TO3Yat0llaUT2drMpXNV
ySt9tpN4N8nrjoI5y/LtE8sbdrfiuWHAkXuyPgmeOiLiw+eWJ1yZ7BP6F5jKOAV69pIr17krYGnm
7RyHR0va5gf203joGoO0d6ffBTI9F5JPdHI2zTAhBop02y1EGtNMTM5WXZeD9N7FDwGrv5Y+jjnX
B8RgSF1Quvi+b5aXq2vDuz3NB/w96XIwMzCgNyTWZrVNeKf+voCZ8F7A7pCsFpBCdv8NPFj4YlVg
xliixkT0Iatr/Fw8u3r42knJ9CCkb4CIp/WSS0j79eYA07nwp8mgwKEaYd8X01v6bTKvMmNyUCTf
geQQJSuwDKiPL9KyEippxdfSfTzgnZGcsGrvN86mxQUSJWe+Ul3Ic0p2r9lC6Nx7tcU71nJCJ4+h
+rOGUwInLpYoUUejHbIChjaFzj38O/LE6YMe/7TY6Y8YHIu3T6qqZHYZnQysoH44ti6BmpGdu5xL
QFzjDzUHkiV1RVIRFtaCbgoEblhLGTmPUwKQlV1K+LzBKnQ90YhsmI3bfiA2LIuGQXATtjhRhntT
DHQxgH+OvUuSxgvSMVMVzbPEy/UiJL99in7rD4l+yRTahn84yVmjq3RVadcVISxD0MrRB/nrMRuv
VpjBKqqXsoKy07y8ZPii72BLJou08dsGUv2HJQjx6kw3xjsTGtrcMJpzVa3lQR4djeZZ5nGBH/ZT
4sQXCHhASOMPI52hLitdqNIl1wNfq48uApVK/0ZWgCcxmGTCXYm0XPNDPKeRXIDzGmomwqtQnHCW
pGE0m+1wi4XmXJ6nj6HJi5aSLX3RqKebcL+GL+2IWQrTFztqPgzJbqGybqEaTRkejVRmA8HJpJwB
qf5IlFlna9l4rm/ZPDw9lsnaAZuwnLbs3QnlJ3r4XQyVwnDuXFNiclHxCVCd4mqqBfPbUjFFim5j
D8zI8oqo/xr07W6/u6EqPOns98LV2kU713CJ0NJjlqi7n8z7xRM5gfkNaFi8Qacbtp3/d5kQjPCW
IbchmDNI2VCGZfw6oqDy0ww0zInZBiQaUY1nKz23UaTjnibnCSw8S6KQjywjkKsDgzSzE5rf8qgM
vVU2TkHAy65iP8y8wEfi8uh2HOYZH2wau9MmoTYYLtRLXYIhAsFMw0aQxE4uVBXRAm1onxN0JNt8
fsBH+VQK69ovWYXOJSE4aO/YtUc8dt7AyD+l4R4EJoUH7A5zIHLXtuOOgOWriv5DdnUoQiW6zUKd
7ouHOhykyqqaH33Djt0NGHI4EhYv0UUHEQwZTL1UxrqS2lHHvvaMn32epCq/dQUuh88XcJ+UPO40
+QaSugcn3KsyobhVxlaM5XqVLzECwdfID+E0V5vTq0vtvpcFkRH6ZmEBLB91m4N00+aHhT/zLoqG
DlYwVXRcwHScrq20Z6SeBN87wmZS3pHYl4Le3gFG1h4c97GUlQToAgHuPGeX/I0+putl14sN7p9Z
SvrUxa6AXivFAv9NCnCVRsPTZWlTB9RHRYjbe5nyq0OogmvePn+Q9mtD82ANjJfxR64fJtBZEwSC
SnRT+L5DYFiZrLBEXJ9ZxBAsMig6RXAJkt6UTJlvcw8//E8Lst5MumRIPbyIdNUeVck7nUIi4ZkS
jvsE0yVWKcnH/UuqN4KEYyjaMwLgawFMzF0rYR+aUkBIMh3xpKdEqGT2fASzKsnSzCgWh6cLb6k9
bqBra6UirYHvPYJmms11TdiBeXZAnxJ8sl2BGA1M8/p9aSZHCwnjBa6a3MsO77cNPWyHppl57In5
dcYKLogJqTrYqXG4yGXaMKu717x8VAK9arD0yDgEe9GOuisG1R7SSbUx5ViNvC/1JziTb0zVMTdC
u6I220Xumi8p7l208mAmStBbyhJleNRFh6toN4NZz1x2wiKAiqshdmtF7kav1uz17Ct4iDTZeg9C
H1qGrQpHBqBDRBZblt5XS2WjpZ1aF7TwlCaUi+oQ9wuA2Ge522+slzhFVqF/AEZo0IrEIyj2Q3Q/
Frg8cngMl4jwKGwIDeb/76BP1I5IXU3EjhxNhIXa5BSQtCnpznPEn+W1BTEevjyWWbi2PH8NymvI
86e8DJQtzRYnO9QihWEIrmwrob3bAL29k5J4571xzcrodSCyLUzFQKIYe9NBSEw6napQPY2T3VrG
+C/SHcDqseaZtoyTPGXgTu5YrR4M83aH7OTQubnkzha7agG+lL9KmakAT/+J0nKe6xMpJEEsWcfx
9Y3APMqyy2NrXvvYXJ8Zt4FfbRGFfv2kvvqFSV+9n89iMon5tAgb9dpiA1HtspWcWkIbXPWAm3g/
alZFy3+WtDjAamDnK063WBtTVQqNfrxW7IyGRK0ZhG0guFLQYHIhAmyuFmH2cuT3nv5mufCw98aw
j3q8JNnHssWsS/dpvJi9OStzUauBTwKwmhWRMBHhK3BG/+c7SLAKrMHbow59NCblLhxvo8v6JzNK
76ECcdn/lPLGvosWO916wg+WOuBZs8aCM3xLF11hJgxXchmZTkBm57a5/YqhddtjIXE26zI5xDne
nJwx/j8FjB3r1pioCwqF0R4+sYCXFSIji+3rJdYBGO1/HCAOhjKMZyHBxrKbWgsJOGr9xnX7aCNw
DYJCPt5dQWC0Vk8R5uXB4ItNqbL5p8nQt5Tb5lXaFPcOYLzhGhky7P10Dm599CqcfOrPLP8mxF2u
R0FO70c/Y25wovKP/EGCBR7G13/cBKek6getL4dbsOoqBaR2ZggStEYWPO0WHQQLRAIMC3Ql7b2N
5eZ3spwb2pm/aQqIF8sni/yGwxGCXt0qotj08MEFy3RQfbLjgJxSL0ZQa+saRcl5Ucbfq0OF/l7x
Up7IOP5zNKuqIjY/WhEGyrPPY8vxPoSTQcjqvo1xfe1gQTm7CfGMADS9j9+3AlsHZSu5mVAVmS4O
3agxRYvTYteVeZzaygwu8Izang04dOYlYNdHpiUNjtfTeC/bOnJG5pmkIlR0K8z7o1EJU7RizL1Q
OoylY1T16lEoOaveio+q7PeTl9wBJkDMw5aRvqAEjdsLGRmrq/iD/1egCV1VC9kdq4i6Oaedz0Pe
rw2lPdlMgLKzL+XHbo9Qbz8UPglGlECd0dEOC+eo8v+FakmIKLh/IefAQulvVD59LOcffCCsrtFZ
MGmtbUgBsetbLnCgzqGMIFoEj7i15XQctCuifNNx0QfR+U4OAmXNgJ6rSfWVirnAcU2oYgPnMZ1u
CbIiv3HbQN6EBs6uGtzk0O5r8DSKpfz3CEapQcVWYqgJhEAaaxlgZfqQ8LpSuMVnD7YQtKbAMSEK
iQT59G5M2C5ZvfPo+nb2krXICA3IlALNBAUXz8LEX7tvAPQfsP/zmxIBo5/Gc85ADYT5tnXrBazt
eeWSFfOiDQnwDW/t/l2rW3ijgorYVkLhn9LensikXXtoIIJ/74jTAO5NkNThzKiLJSW3pIX4/OVo
UB9GA8M4x9GlGUcMnLkx/WN3DmSj8FcTnbIDE/hStvPSBmStBUvEN+JxxQ0Hw6iVBoAX3hV4IBxd
wIemxdrx+wq52JPB4OaC8A5e/sPCAB+qpg5mk7p7wfOSJoqXBZ9/w+j1U9X/RAS+02NvNB+t0q/t
JfckHFdAyz3rq04Ea5AfjckFNQS3S3V1pJmbPRt+w+HuL58q577PsPse/eF1SUzpV2H8O5HA7QJ/
MVJRf2CIegN3kl/j0jgpgtUV2RA1PY6bvgO9W12JgbdgC4Te4UIoYFJ7OGO5sNrVFsefiDCdW9n2
4p2lcPNkPI3Q3xuyYtBxJk4UCDTxQGj9OFDFeTXLzi/j7iHJ/GRlh2H9O3w8AyuOkzR/BLstlF87
+SpFARRpBFoNPvJIIfgv1/UOCBA4wSG/vTOsQed57Qv8ehD1Tq24CAEO8XEEW6V4DLyJUNOdY4v/
rT1O577btqC8PQbkKlofNO+cGnLoJLspssYaxvuNLP8p+oCPmRrzVgSttqYFNEiWplHBW5eiZAbM
XKsZdrcPYtS5CvistjEntbwi6XMyx/uymexIqlV3MEE5Uogvp/vrDvX2Upe5L5nXwKgik7qc6huW
ZRj68UWynoiCvlhcL/c0lcgHKquaru2FI43JCENy+w2iWRS96IQNhGAlC2xeoaU5yPJu4Dgg5aIR
8/gu5pJ2DmoKviP7DQaKBixKL2/xjOHOwYsa8h+xfelPwFAiLm+NVthcnAmfjm60oFqrsjl4s6H+
ODrllQZGAgWPoPwUO05YVMlC9fd7F6/SGbEl2KgQ+Zql7TYZkpo27fu0WeKtNN6E5X23TLMz8u+g
AAeQ4ewmSIaGSIMPb2N+ZJN4iHEKoWvlcI7K0xyOmI3wSJGEtmeXQFl7w0x3HboNTKwh63ldExlS
qG0o0LQI4P4XXQog5ScqbzGw1ujvGaovKaUR27Qa8Bawh2VO68JoC+grhUGILPwrO02Pvhozy8vO
cqNXiTOb5vMsmL2/IiU523Xc0en+OXuNM+pMpjEaWbl9BTXV+DY31DzJiMJCe3Minl9KSP5o+qtC
gl5pCwOC0WQjMP+323JIglBXcINnhGHQk9OsZhwXivTHt6WTp3CHbZrkl+xntPHvIwVPzRP7Rs7X
08mXiDcb2/Mv/Ne5+ELBwPydpdEEbVYjnxSQSeLkLWWvfvIE8Z99OQ8rkNObuxFHsUiaRnJl2vdT
2OiJKm1EBF/0PyoWbC8tJQbepf6iAiwB0YpHQ7emESeTu5n5W1Wj7nwvF4E+4CIvEie2x56xCwV0
sniI15PTL3t9fsCx+99JZoVUMWK2NgOQhrPXoO5SAkZfJWl+QCSOXG7DVeNtRRshuPdsKEOGwvyc
jfLSskm5JV1PKNKM3NwuL4G52fwNTU0HOEnLGyoX+NbStW/X36IAdn9rTAMSLXvxQ9OXRCCofmHi
QhZyQr0nzWdhxrrlmklUfQ+BaACcdb60iS15ZC1Yuxwwm/mp3csLI0kuSKZTACrX0wUEiyFSCNsD
bKf+HDNDXfK91sHlVtVfkCQpch8S+ng7AV3mS5/aKQiAJDoqelqoz1PJeBUHtNM6Let/Nld58z3C
dN0JJJmRas2HmK38egCcKupymYLzTEVSbxP1hOkorB58MDK+UEG5aX4OjD6EsORhqCDBCaDNGPr8
ctmK0miSFp1cjSGy/j2+Io+avIslH0bvDP67IDFXxl3SjzX/PBieI4zlYfnSl8bxBjcNPIOYlMsF
6uvymMYucYSDG67POeV2peGRPMi+mJvbjsB1Rq7S8qCvfdegtWk/cnSvfUq7afrSJNqsrga+jFif
e4REXRu/b4YB1l2lRrhtOmX9wrRftg5cDFKhzNA4wO2RHDBG346216IG2rw+yLoYEopKnO3xrUM8
DuiHhTBOzlIewXNeLwD95yC17iCcE7GUErPT5jfmrujVhSGpY6qOFufKQH6pMUqNTL1gpPBXXwQs
zRlac0aEcoOhSMc8WEIHkhQzOan0TsZmKZNjQKy0m4U1kcx9Bo/oMgaORO7ljIzZkdake4b4QMgA
z8FYrj9341GeagtKv0auV1ksstDW6Tj4SZX6YOmMnCsZHOnFfd8B/qJ9ptRDLh1jXWSl7LealF3I
uf7zpl4oc7t+PJsCSRyQwXi6cfDhiHZtZ2qAnr7/olWfssNFL/OTJ4adj9vthr1Rq98deXDsyH9r
7XbHktJleFOTAgRGMiIhENpki4CLlPb5ms518d73bSTiErBTDHEZIi8nLuLdl3PlCdjn0rde9hMR
dyNU8M1tl9fpRsL07VvIzLTb0zbLfIbd7kf0r80bg/5lz8DgVIO1rM1/PrSTugl7GXsZJrMVQQK0
OFSCDqrBaxh00re36uw70CM8CJ+B6EUNmWxBuipZzKmsGzt2xNOHIKmowQ6eNiqiPc2KBzLEjZOD
+OAf97r4z4FH2FZ5XvsX1XB3KLa0baVHE12nBfqZo85O7mUNj5OEoZC7XMo5NijgMWzHuTfVSI2S
Py1qWntw1O1aCPoBQkh/czwnsE7fdS9FeIcboXUvBWOFwnLh+4WqpJdxWc63ew4Nc2yiUwpu3t5j
Mi0fP5/fetx+659uJYZL9vKP51xiuR9a6Vpzbc6154CufWMVZLsf/Tzq72oEAJQ0PFQ71GTZb4BX
ZT0bQncEu/7r6AzJvu95fH31E2JgJS8HhoWGOvD5T6f4qtJPbbbU0cE1S3gISS/bcMZYhv2bPLy4
kMqGLk+1bBlEToSQqOwxGciIILk8aLe66ScbArBuHmxW0gTt8ysfiukQoKA+PMUIE7WaQpeyCYDN
OAXyGTEtrk7cpMaUeRKhwPHpIANdiE4kP4cPEz1Dp+Y/K9Kq+WLzYxj9ewq1vBolCuumU7Qk1Avg
J+FslZDttJJjtRHykjPKWXEPb+GkQpFjZMKQrhyA8ZOzc2xqOKy7o7aivgBTTiF2OL5Uvykl6BTQ
ZOuTC8VYfniJ+oN7aZ0cpqsoYLA0XNuPj+qZPa0vVx3c/24IrVDNzve7/o6XeKxlhQ5EdksY4kns
2WaOpW0g1KXGR2hVCPpvlVyiOZmmfvVvnUV/ci3cS6vdtVNUU/2LJTo+ztU4vb9R15I0xM78ydQg
qAyi1xt2TNmrJa7r/HweWa8RYzGw0mFeFy2FixomgSNUV3dpUWFzMiqWbEFPSLkBrhYswMt77BuK
t/MffqlTzsV3ujKUI3ZjLXBoBy2OuUcyOlZ1ztAXYq/xTMOi5LXOWCgccSMLZ7sDtSPSbKa3j8Q5
d5drOk1pZjXCZVknqHWDudoJb4d4crEzPGeHYKQlMldZ1GYjOOuYBQGw10G5fTUrmpScUDtlupjm
nADreKFDqXDkwbt5K8ILCxxXvv+DsyIBu10pPd1r+j/x+vyyDjKJV9ibcMwGyBM1BiGo3U+GyGw2
3lMy0goFnVtHvVWSQ7FgHLTvImYXTkkWpHqp4ftDWzdMpwOCmwx3zaUveOLpSpZczRLrlSrr6O5y
L+tCp6pEpjh2R4LCYfqsF07jfFFNabyPBhjZRyojbwqhcCtN8JEKopxkPWsMdVWsi0GOKZPYcJra
1LKNY/Ty/o+0xKYfwAxdhLZHNg30I8yHvSW1csxlZp7Q+8rfehSOQLbHPDxcgLdg4QKFmOuEL+0C
H7GzjxdOEdgnT3EUWX8u4GJ0ccHrQiylzHReruAUJTWfix9Rift2HnHdolTNSoANNMugEsqQ6MAF
yX8MhoHEkisUl4AuQSKjpFWXAoRpatvrHXiwXW+7/WnMS9e3qHUpt+NluRB2QLp7HqZOlu8GPuja
MRJZ2ct7w+nN31uXYvjb5QL/oOt9HSU3Zpblp3pnv9FDu8NuUrVFas2Yt+5VZZIub7dWIJN+ctrR
1+gjAl8TdDXrnHv8cAo4X6xUUZvwmTA7kxvqXaADxflKSIoymta+wQZhLV17FpTq9cNFWZ7TT8w9
U3URUr2GTTS9ReC0YDuvm5MiObGWy87nequJvQPPRYviYW3IF4zNGqKByeRFFDe7lRptDAlTldKz
5yPyNLVjYqNqXW+7qlWuA+5O+3evLsAootRSTYOMFluBsZUf70HgbaSQnjz54q/a8niOJFASlwU2
V915m16Pere2XmCwMhgD9yAPKMpa3icIb1WNIU/kMx0itdt4JUifbzf0Z2brcXI2wukqQKfaNg7y
cW2ooZEhu/Qz8NQPW9IoOCGEsoSTSRx0Px4f92BbvcxBcXKrnlFAHXYsbuze3h6uGaj2asr7ZsQw
xBkadqNkRJ0wSkQdCWLTc7H8ZHp5ZHb5U4oXmMHhwQOhFfjF/XHLF1AA/8CH7Nb26jyQSbmM4DPl
f5eOzz4BWXVYVSHaJK8a/GxU9WJKs4mJZwAnlwGR1FVPjLj1IH2zw6mVi+y1OSML4sORWv5s/TL/
irHpQjfYBGL0CjVDDh1QvhHawA66IY4O1jZ1B++GHGCULsIk0MxL2weEvkQ480I07vZgTUiKLkJW
jRKVXivZazCyiziFzxiSqauaYKRZPdvKcCBaX3jjzPsN2kjfmKUeYSsAUxODHeLH6UHN/Q2kfQSH
7xgoUzzRU0J1FLDMDI6gGlwaNilXNg7RVJzL9laJ/T0tOrWCfkGV968zA584yUgnthyEh/mdkxD/
PdiVX1NaklsyF/gTa2DF7fJKLIejRZUTqeeUZgK3ayVCyjyE1EWKJMo3PcRVuRYmIdTdTwX65eS5
tS2N+dR0Wgqd2lOfKhhOKDTn2v3uhrD5E26zdsvGrjGXvFxEqz5iyzlcagyXyD/rNHU3Ta8vEsS2
5JJZcnxVnSN9azEINSLVnA2e9eycynoqQKkUZS8jJqC26aGuSqX6+3fLrg9J6zaNrF2ZYeVudE/y
UfQsmSAOXkS5WYzPie1kGUTZI3Pxmmg554WT2aZwM5ICikQ5iDssCtTQuh3U3uulQbceoTuTKLK+
WXsTn9VXakW/Zl5uK4HY7N3SFF5iBjcn0MFWHZyuwLPVIN7U2Ks/VHROdKKZW/CFFqkQluP0jU1O
LZ6Lg5v8FJ6+MAfIbe+7dLdjeB5zjxc9dBifzzSp45Vsp25urAihUYD+RRFAtQP/yY02Pc4DgPcS
Hm/BRMuyr4etIztjGAoIx/Z0TMSdRDFZXi5lTzLg6tb4kVnf/bo5QPL7h2x+2UgNznzxXd/sfCOn
tP4LTRlnT4miPuUsWSziEl70rucNXzuVKguhX3I17V+82qVr1k1aZlLi5Y+e7Ok7zm7fmUb63cHp
VoR/DB09f5cLr+6hX1yBhEqmUekvF5MIcH/jDGobvnUW8x8taY2hTkOHdgi25MIOi54lKNbPQ5FN
egI28pHwhK8OfQ0NtHb0liSd6EcNKQGfrzkzTYDSpAQk+n/h++/uFM9YPqZ48pP/5YE6vQqVyQWj
t0b/271tD4XEvcq7ctDkd7RtR0sKyzKoZX0xk4blqztpo7F+djAEGBQjWFlh1BuRrNxIW2zBrDjk
uL+2Pf/y1ntPAvxlaMjwuQZ85Fm8WH74yXGOrA+n0+Co46yHJOlJ+6AUijWOr4sL0Fk84/Kl/5SB
mfkBUUBBoEa98Vt4XGztOwhBbW1x2FynCwgjqjq7C0nPRI7moeJ8k7Bz86F1geHkfaAvLXSSyi6d
A4tStvv5yY2YMBCm1/XPaN7Wit8H1VXNWBlypULGcgewB0qR0hkDYomMGH0SrYVavySFf3v+nDQy
QhyW24AxAwSwSxaTl6x3ZBRcwbpIkvM2yvhWV2UOuTrTV7qWO3eqHFi4JeWVORA0CE4y0/71YR3n
XVZ0oeo+DFUxut/mYbrrY7X/Q/1xzsCKmgWqo3s1VhZhafPSxxoOwtu7LXLQ4WbTbG4/iIgWcl1t
tVFKCVtWmwrhr7UzieV/lX9FtJSHKCazXbSwAx7x1ZB7KOAv9l9YYrHI6G5g2WOdcR7y8zEE7Tw6
iuq8Ve9F/EsToL93zzBszk10/phuz26D4GDC5C0oSQUuCMjOuZehdNI9+iElTgpcs/TCkv0hCAyK
VfEll6fqkBPhuHfVIReN0l3MGsSmaTrcElc6juSKX8M6LLtuZpSjUi0jrDzPmDdreszyUsCeP4oz
T176upSqyvGGLXQmrpim449yCvc3gl57n6NSw9ryHdTeXSzbZZVWXl3W3xjhALoU+Bl5ma3OHeeg
ZR3JpYbzjOm/jIDNdoa0+fYoUoUaF2BLr7yy6Vg2m59awvv6SNGQSWI3D1sd6zZGhuSiGoAcWfVQ
9lL/R6QMD1Hll5SgaZ8bNsa464XF4uwSRxus2vfZvK6lhXOYDwVqAkLTXpgWW75VFwRRSeITsVpL
m48pYZ1TUhNYvjgxpqQ7b6qaf/O10rf0tLwk9anRQ+6mu2HQtwOpM5hDbtde1LXNITnexeHvjZa7
RludkQztIAxHx8rUBApUmwxP+CgL0KAWvNesDa6hJWQQGXYMy4AV1auqrXlGxASHX6X48z9RCysZ
4VSecBoKEwngrEBZJXu3PJapozsKnaWNFVPgydztZCNM5/cmGXuSb6aE6mFIfEuBceNGF8Rt21X3
A/LLNcoiUE9LESeJpP9QetfeL19lFQPWFllBNOhfKxUbPAUi5B9EiaGNhybms2LWdBxqw9LVrbp7
2ROQUsv+t36cncDtWShsrGjq68/v/cV9F6nSYm/Kx0O2gQbQjazN7xxi+9P9DqCQQcb91aLiB8cU
u2VWSR6wZNE4vmfi5DVxpRv4u87LbEvZiIAqRR7xr1FbkX5BHzGkZGpjsKJNnaum5JjcFsAspxjF
heH/Jhm02bWywzx3+mKDeWrDrhPQudyaEmXw7SEGrgf8or34eNS8VmZMZg0+Zu/jGhFgtfUXFtzu
5X81Pmr3Ny10YmLh+8tYrlZKfU+7fjEoMZIj6lzMDL48RejtafN0XtgHTq009wWPeEXMsXP01w/8
VRxp7XaPAjAnxxmEwSN6P0p+xCdhHY9QNKwM8vZrS5ZUe4uOEPeMMwTQQa38dFy3MIdH25O+kcBj
0CQx9nLMPi87A1yue1WlO10OoUBWUEQChA4ewuRoup0VrBwPHP/9wv+/lOKIk3+rFHiL8MLjYhxw
RdetQzfRG8GZ+tZhenkK7E7SWZqNmIkIfzI87/nIwq2L+aOmozqxm0jVpV8XgyhcqEJeMHvxNRzA
cVXpXvIMsCZYbwsk6aC+ooPRgXc0VkGd6ojJV0kWTwIBvCSl5HOrSAGl9+me6wgRxodsEfLy1hmK
1MbuRqPOfc1Ta8qVWDy/d05OyCZtS26y86YuFSZ2UbxOrG5GhmJdtNO+1pGDvMkKIifqgWKhrMFn
3TiMprvNJeRhKshKglsbLjFNJ1RcIEQeVMh/HP3ml9ZjFanjUqp3hqWZvNqUu6yZJQRZ/1MiaXM+
OnO0UTKOYANeRBMRz3Vfl7nVPZVL/8x/BG87tl4MIBSvDrNN1a0zHeV/DPArCQnQ00iGmtXLbXnV
chSUTGnPd/uxKG/ngJEMun7EJZ744ME7pk9Lb0lVHgNLRVbasS3ND/V2ttF9GG8yBeqaSX73bJjo
XOcDmlOdWdctPr1dbjAWm5cGKm/9Qjmax3IFZfmPRmFP76lMemwV1IgTentqjjc5rtCnHUj+MAcd
7Itn/K7UPrq2K/ktTOJ2FzOrITkRk5I/JaJqpWZBVFDztaDUYRcycVP3aEv0O4N+ydOFrIfr8MlU
QvjFYwE9GffP2Mkoz+rwlP3oVSb8788Jh0wlVczGADNxSTp4Etv14lUcyyvxU69qFkmlNSTgeyKb
FhJby8N2SMPRit/S7MP70Lnpipe8hqs9+GOqFfrZfBVsd21tScIb8eQKlN36oUUAUgHoEMareYd2
nhD9+ymUDA8vEGnkvUcBm0bGkLbqJtCmmJRYoADxYYRnigHMDMRqQX4cQC3WgDnDDk4uSO8+1YqB
Za4pYQ8QV/ud81iNbspSunU5pYj/MY0Bw/umbQ7hhob96mJhMArZq400cLGjKLxvnEnj2jqInv6o
lmvfqVaQbX+27svQ3xqI3IMVHdBOzqe/kj1jiZINprCLmSsWO6kg/UJZHEUtIkqqaGUir/n+L49Q
zmzwy4E9Tu6iriJw/87CKVM0Y4u8SF0zg3W3bETD0zjrF5rfvaOmxZA96OcIVH1QJSZ1kQcyUOIB
4R44Z+RP5tsgoE8cNcEMBFliIfjK9plt74THj/xybz6H+ts2HJQkH3eV5+4u5OfEcTaPdXTtj3bl
G2EyFedZEHavOjRtftIl+A5t/xFepZABycZuxjoz9uFdMYmrNyeuekag+g8GmAxVwzSjAh4nHiRK
kp/7xcU8S0OTgFpYZfe9eNDGxCdzAuY4ugiaQR3B6abH3sIswDhQmj34j9mFvwCSz+XUiXb8S+xa
I8+44qywDfo45kaTacUnNt5VVApRZSpozX+rmksGzD3oM2Vegod702RXLzYcsjEYpDJQhgNCQ+78
YvC63hu6RiuVFVDzoZX8lCiaZuKPkS/uRn7I9id5jM74qRVAtPGYGFfFRsfSuTJr6Viqfw6EbSw1
CY6VQyroT+UWnF/P7CJOMlT247ocWmjE+c9KcDpobQDpFhWlXfVc1IGV7XFp89g4sMWfbgfHBcJH
uFt9a9FI8F+T8ueATQqcD2WbkU/Xbk84D3kbUkEbFB3r2lRk9pSdjOuCELiKX7qCH/QiOrVFpU+g
mOskxN8dJIYP9fzPvYM7TlOvcn9oEdfbiJWWgubk/IC4tDCoEWPu5n1JGoVboMwR1kkPbpziZGbH
jQSZbnmuB7ANypL4gQg8U736zkkb4K3BhoT8KzDlw8jqGe7Qo2Q/xHqyoDzmwqRvRu9O+L4W5Tmx
vKxjXOF5iHiPiEPcU99r9aVbQ0xVKuVc6MKo1XhQ0WDBbGTZVPKSqMRo9iyrdoDQ8zm+3QIQ3bGT
uYx4Dn9p1XPFVxJtgGICZXQ2H4XmOrUi+zcU4QId+VhShXoSG0r3fMBb22A1PK6BaEP1se+ynJqT
/UeriT2pHU7Ba03hVJW7f5MEhWFevqa/kP0s8A70AV6uJsy2Cbeys+2delB06e4nGtLO83vylXJE
dTfU4/IFxESwqFQ5YTpxNhd6QU2AR44lwhsaH+ccLG2PO3Hmy6gQX05mXLGyJ0wA/g4WMlPYoqFp
/PVqUBIQh4norrJfSv1WduPvRfqwZD/e2wNEoI85zmDOEU4LOfiia5S3mj1wezmB+BZz90ZXReE6
qH1tl6yNIeoIG/tF5VJM+70OrtutvJ+UNNxV3Tz130+dxJRHatjH1ZxdQw0ZOovk+Ey00iqupAAc
K5Vy1lxyHrvQTOf8QsOuyLgPNJekJYGcROwZv1kzu0eZjowTo+VoCPwe9oDI+s3VnreMDg/9yYr8
FUnTSN5eYH6haK3JD3/E8HLcpPKSynjYT5EomcBD344MA6XCIBmWTN8fB8Vge+AnwUGSOtMK9Ihq
heo4QDh86wSVPk7xLNTt+HjAsF/hfFz2oj89ffneNRNWGPAsAz9TW96+/a6xhsYSIuBxexSNGU1x
mX45appNE43nMmdRZXgd80FknofqGweaOjVBMxUH0FvtmMF0K/YHWrHOka3BIQsyyO9yXV/S1DYV
tnPCHcT7oT2gk1yi8j7Fllu+E8+cQyN2OrjHx9RpPIZb+3+Y0Re9gQA1Xag0kT/924sIYlsOtA01
XbYBHcQ3HxiAMRexL1t/mEyqE33gwXbVVBPkSFgnH4ydBMq77BW9VunY4dgDJn0L0DBkOL0PaanC
IgqgOjdUSheOFMseeac2JtOVhWGGvibqKEAtSX4CFxPMk0cG9MhvLRSw1E3LCpciQD3kTdbz6t6W
2OEcwXKG8qYxXgRoV0dS6t3UNDRsYt8/BLrg5rAo0rGTro0uUAawuDgGCzgXqG9dpQ8lrlwO1xLr
QrEPKaG0RaxTZvDjf8qpgQBZyVD4EdYEai1/d9h+19lJX3YgS3SHwb0WRjHfQu57ZgOF51GKXgNG
oNKO5zSu5fDdA1SiBBKo8t4XnTlMEpDoN5izcrntfwqtxZUN0QUn3MDEBEXKmAV9WziYAvnBUz6r
Xf5DsWp6Dtl6YuZvhWXT9h2Heyfysg5YXF1nIVWAF1WcC2jf+LwCkiUwwglvC1PV4G3SI1QHfXf9
QD69yyL9cw4ZEzMeOahG2FJPic13/cbd1tSx+l0VuOmm8ZgAsMAtM4PYzx7ooI/QTcOYQeSPHy9e
dfUmBNGh7n/wnwugkVGxWTjF725eLJEEDj2RzcPOksYZvbfftk07vS8wR3r5nzeWolPfVAwxptXK
ahpMm+HeWMTMmMdClS48hzvVz/AZclG+LwdPRvAlwu0NP3UNrYQwdg2eP2oKjyOiHkCc+vO6Xy+2
aXedYwlxfrrZE25U+VfjdHuOMsEnAcd/C08EBgZoAXBcV/uefaBaVugPikDGhUtODpPQTlf6ZrMk
Yg/6S9sDmgk5htOh+D28KNGGwPlh73ER/TJd/IKoHMCRQC+q7bS3NqvnkQplgP5RkmTolvlFEKYw
eOYyvbyCqay7mqaNzFWW2kCgUmHlJdIM/YHs6gv+I8Y9jIEBsfqk1vKBx6L9ajYg8NyrFEkRQWEO
280Wt+NdVN85DNa1x42vHZ+sc3bxQfR+3NyKS9CmnHNyIMjyLBl3D1CkWdyzn1rCITBRKvV4BMDt
d5z1DaARfo3ZSKUhcNJSx/tyfY9CL3QPx6E4bs/s6UEvbw96lOyqgO8J6dg4hxU1ANK5ydvmcywT
MiMshCya3c77pedGNjqyuO6NuQCkZEnGk+q8UUpdsGyCkz0deE+lcTpFKxcJvy6tIaIwOlTIED1f
o4fZujqcUx9CbJa+MK+uNNnby60mtF9N8d5NUWGi5ZpWfEgJ1lp3bzgNXvynaYj6hblRnd+MAVCC
Kp+lxkPHD5NTa+e4eBtSb+vop8iMlX8+i5dHCzH1/OPHHn6ezj/zd2YAvXfWlcCA/rOjrNmspJz2
Bgq2ITM4Iy4oEmn7G2DJYjPdaKtW2Db8/iwChXlNQM1BMFjSFLbEWF3WCiIeVrQV5x0XT+oLUJBV
KrccifbTor6FXGSlZ/pKEFVfvdcPBVhJQIljC+fl4AQRwAE+hEKmFvA22XYXBaCRaVAsWEAbBIi0
mivJVkc333dSoS7bVe5O6YhK5W/LYq1X//PQz/XcVvYQor67ZsGuvm4rYoj5egWyKujARY8dR13x
EJb4AGHQwVH63X1FtXz8GayLoZxtalaUyhI5sM1dwnnMAa/0HsIjylyDYij0rKEflLVpJipEC8g1
XJ9yZNLXIdfMWcxqXY9HG819Ur0whjiXoZ3n7XUKCu48OkRA4pXl4P52kaVDdCsMSIhIt5GVbct/
In9pFQNQDb9IYI7UT29rCiwsxcEx5BIcapQbE02WYxMHwW6nU+ml2LS/rPbSXjzo9M7dbNEKi+9U
Xsi8RClIAxN92Cuwv4ngUxacW5gbKQtIEnK+FiAk8fy2633+2J3kXLQbiDl2bgW4Vjl/cpDoIise
hvBqyPlsyLnhaV7RseDoEv7IeobsOw2xA9PG2+s4GcRjzms5e3GAFZb05gWvo9KMF3l5dfqJ/kCG
Jg+ecpMB66KKDVyX3xXOYZW7AesNsX9pwKXk3hq7w1V9H0LB7Wx4PkyczmCsJU6ybCI+yLF9x3n6
um4HB3eJaUV7IUTJinYQ/7YaC/61PjAm6jhxzAfC52KsvM+4opFEikn4ehskv/EuL3w9jx3htPKr
iaIBHqMw4lkgE5um8wkmIywplfT5a+ggyWSA00Jpg238yE3OQCJ0/13tI56LzFjeZS8rvcCDEfYM
NyHTTn0rrhP0kkU5V1Tfjls3gmC0feh+Ga2P3kTX/8PQ5SJXyfbbbhwyIhPveNwFVx9qPy/8u/MP
wo+LxQeL05P82Xdql2c7NheDG519YacvdgL3tGV4Q4pU6tS4DVUwXKJJ+/r09893otW3mXIi1coA
mKvGw31f7vvRrmWn8FYztDw/ncb4iWmS9XazqLAS0NYcTb9vmJV+wUHqy1aVk2CfXZSy6LmBLauO
348RBHwocHE+PIUvUCu04ixQENueJayEWfl1Y6p3AAt2pPBzE712jvec/5nOLPs/FvXrVOBOqg6z
1NH+UY1TdLsGKlqBpPoLvPPHq3R7BcfTyV4cOTa37BAYIexgweC8lr/VAwl4wSlQlBZC7DtkDkmI
gfxnz5UAQX0m2cU2nUOPvgwfncA6B8E8Fc/GyU70gGIGTSj3avsXlug+qWB5qyy0KNtJcOQpVIk+
8/XK/bhJdQaXVVjT19ZLhDQN5ZGHgKMhgseAurq0v9TWVuL4DRMCts/o+CmBBLs+UJCSu4yVooKj
c7qrzpti2ofI69HDCd8UQepHBreJRVya7z3FekOK7wKBPzFerVAldzA+w4oKoCS8T8RWhsjcv4z6
dmLXiNuDe8IDg+tSW+Qlt+dWLSkDmSTWIk3mv/7Gbeu8sdWWghq+89YLIVnsIZBbWTTH7GDTNqWU
lUB84QTnqJtuoBszn4O4QoZ4sRU57XP/CkQwMpXe4h8fFUHOVk4GpqEI3BJM8A/JXnN7fO+BlLRw
IMpaMsw0+cRuYIBec0R8nYczspx3nxgEskhI+fXgb9TkyrS8LVzWJM3i/uJ/EGlB5MuLvvW/PrdV
yHSlpm6xlVpnms6U16QMOpE6R+MXPZlQHjcLqQ3b0UL6zAp1LvLKuDNdtvVLHFPWedMaABfrDXPq
9cgsKe7RTrncyREKOwuG7qSd0bNTo3pJ6Tt30h1wGnLGIAJ8Wfd1/LzREzJF20c1ufTaLpX02vBg
LrfYv91JNUTAlqWRIP66B8gz9zVBXPCZoN8lMr1ooPiNx7lLncwkvxfHjHY5PrKqYkRsoDuCBu2e
yp+ZOZTxO5y50lh3wpoei5iT0+s+AvSXMqHOZkcOmswVf5PrfwipnkbGBryKzdBkwweVa13jN068
xjRRE56zUj69E5NEuu+iNgLYkC2Uw5UdMUf6GuO5OYA8Z8z31dY8Wr0PFZxD9WqCSt7lcp4ANpiH
RP5E7LtvRK/inysxjed/vsVATKTTdayiBLTWsQtxmRUqetEkoJwlEjxcbpmndYyNXz3pBuPfZdDD
dlEozRLUBWZzQo2/fjjm6ROimsOaqBGYb8R9mCtNeRzivGuBxtWbjSMh2VbhvoDXkeUfNjQ4Yq1i
2+CuX+WBekIBaH8jyxqpdr4lRyrPf/gXbKHH5gFIrr+i2bdFT9E4rqafYgouugYvg2weJ1Z4OP94
LaCMTddT1emjdmWfDuVJdjyWBfluiO4q3hRJL/x+FZ4dnqsDuo75sPQ/0CTzNk6DimiaoRUW1b2z
3zR6of6tPX/2xvTm+fYRyOSjTm86Q4cVpYRIJWKVykuNkAfRqY9vHEy+dpsTElpteEkYmPCQGKWZ
HAnpbXEUOVh8CudFMMBhr60BHKhRixYqL1lBMSe2X5woY8pr6aZFr/ARK9Q0Bn8OVc1NcCTRJLSw
+cypTj0cDU2Y2c8GmjrxhhDGBbciLcszRlb/qaJqCYXlrJd+opdY+wraHpug+9kLkO6oxgoB+3E6
Nh+XTlZHvACRq+Qe83UNKJlHizdH+nlI4p4YDX/s83IJG4EeQ/FkQcK8UxaJJoJLI2T7nVlqfNJL
PIqckK0ftqjvZIGxlYY7BMF02nc0q/3dUR8d+0EugqmDngjIMe/eXuPjFZ9gD7oS8uWSZZJpgCa3
86K/YQ9CFPki0O7qse1Z7LWl+0/B1/lIBP/3paEDWv7EKS96oE+YtqvpZZI4mdHeQlFu2h4GFibv
38k8Dl5jJA2rMkjUcaknBoxYfE9CIGNv7kocQInPiGzq5Y4DzTyuDYI9hnRgSEOnJPcGbtbec5xA
H8R5+x7AJJbAI5xbXIiKfdEzluBh/NY6eSza0vkZd01XIjBw/TvQzC/JVfkRFMASRBlgyPilGKB6
JDvCHEC6G9ZrVfEGnuVYUQ/e8JuPX70s8rqOhaRStQ6Fl1o7gMr1TBycN/gF9kn2gKEKvyzD7Pyr
GOP0/wzohfu8PcdSFYXFuzBHJs4HXPgwXkwyed2LAUOnx6MaAPfBXnDTvGpn8jcA1qAZv1evWzpM
/SJ9WvDglksBlqXbvCd7mZ/wiTzpQXHfioUoArd/XbEbyevBCpokqDKV1Cfw/UW7jGsuMSQUDlKw
vTCq17UgvNn83IqIISdUQTe/X2vZtxokijmRy0Os8IWFLlkfe2yWAYk2xr5lkzXROhKYeZEAp9BV
Hoap2OoAsSbR++By5wRZNkx47i0sCnrNZp67Iu3ZuBv4nJfFv5TaurlNEUTNahpPnDkNWPzVNNU6
H8sVIXTX3+Ep3bmxp8AcvzTzJm4OjsohpWjHd5Oqx3aG85Q1+14B1eSO7dFyUHn+spxFVNbBP+EP
6p8rxkQkv+suI0EI01N7dcSsAkk7eJYCNMIrWxXNU2gw9WJByyfSM0eX6Y8d7XtoFgThmXYJuq/d
vPhTxkX+hXHlwE09MKmM0kNC4T06osCq48KkHpbKr4jz+t4N9941uSe1JGoOLpGV3Ie7P53xwO9r
cr0b/8bqhaRoQ0L1KvJgDnhJlYlSQFscNXmE/01mRnPsB3/H7OiyqxnrBXeWywYSJADNMaEdPDaQ
cOxnZ+PhjrNhmRY4LYjl+udxn10CMVpgCV/sTKt1EcOcQnOnd2+1KTmpWRcJdmSWjdB7n2TRSb0Y
VKuBDxjNeMBBFVw600OapaSP/quieAJAr59CitXm3b0mYK9PhFpTZraAuZJrNkaRRhFUuIz6pgcJ
rghxuyb0MbRsmvBBoKiDrY4QU8TExdUnAw0MlK8pFn+rQz9tBXf4kiC70upDzSeTRL6yzIcbaWl8
SCpKqaVkc/CiQ35gEaDKBWCZpVZ/rfLtz4kPhte/+B1m0RrvdtU7DO5a6Mxrlr5jq1V8GqZPS4SL
FHH0p91QfFcdxrDSSflqz69hg1Y1PEvo3mrJ1eCC7gmscEay1+T6TWGiQzqETn8WmMUVUrk/TIcE
Y9lqScRShhGTrOJgGm33p6t80Ti/7w6Y2ZFNOs6gk9WOTavZMKkelSwWhXYjbeRvr+58tlh1VUiX
fx4Z56kbXS8z+oa7Li1RylXCfuQvN0qiBNN3UDJsRYxgwCbFdis0vQnaQ/KeyLAWC5tiAvC4EN2D
F51p4exQx89mT1EeLE4B0IXOi3TTdjwGFtA/dBBAsVne6JhlrVPj4LuuI19keyBKCEvEXBNitujX
dkkqd4UQ9p2tFHuBoNmBLNgkC3SGTSEOmYt/YgiBSTc0bMap02FCxiFKZJiSJwJiyrlFHr53Aeqb
oI8ytsvbqr/fRSoBWYcr52NvtUBn4WJXBXXZYxq4xCuyo+qUsh+2jYnCmhBRSHzoad7VhrKgrgNy
cUnhpcZY+T1AvCh9svRFttAKo/62YhI2ntw2KiZFYennl1Uo1p13T60Ki61vgJdr98z80gF+oUTB
VpvI7GOvuui0Z214bCbC508TeuNusyCklNHhTp4Om1raQrpEOssEEyHzINcdUfwrbmzbq+/AZUKn
lYhz/pTWo54i0BYzPoTNnebTsey8krAmosfJxER1IZDDlIs4SvnUA78sJr8eKnS/MHCdQ79BRj8Z
oPuIpsj8mojUCRyIH3EYQtzBHz5Hd4jMKPHqKtWdc5z56rd8Ei7GG2+qIb0yL1QMzoOoVki09FOl
ecfcrwgPvCVu6PD+VKSraeJZwMuwNUXUPmismJfCkJsMyQm22CfPnmt2tBY7apeKkkut1IusegwQ
t0WPMqGluUxOsq/WLZkrkG7otNINFHAqko17SRu2yC45L4F/ud1d2EWow0s7v4zmXhb+nKA4+QOZ
3pqg+eiv3Px6WgJR2nODPRPAasamz22haYBizq5braHnhftCCiNTDE0P7o92+KQ+2jo/ubF8uve9
/q10PhJfi2VK1zcS4BKDvpg2obqu3xyGMJCO/ozwHfJoDI2ppFqSCEKFoJM7cD8nN9CerCYFocdq
5voqBfaN4vKh/hhzlDQzMCn4z9ZV1IOX05rL2cf+/lZe5+az3N9yT4w0GMJ0aB19tIasPNtanSoH
KEbOd/pPnBWjO/m79DLNPANBYwdcIMjOZlTiF0LKiFpa0YBnWExKmzsq1k3JbLPBaqqUNWImKEAk
hEWpB8T11uUgpxoI9zS9c+HHoub6bzKbSdtkpypyuhsmMbcnscmk8+tAhfd6rtwe2LX/gkekp4Ai
NTgz3i8afFiDCtNaW1Pm9dZtV2KHVf8AGxN3FCQy33MfkVRsZdvJgUi3OvWc5/FBmHHUfuDaXCrI
SeR6pUBnhXagrkySilgFEq1cTS6LyvOdYL72oF2TlQig9JuAGryAR9i33w+2SQjt6PF902Q5c3JV
EWl9lrDSaPm228LJ0yKIeduBAtIKVfNoChoGLeObKupYCdL2rYFQSNcnPZzjhLfNvb/wDkXnoI7T
xT0tG9OvDMbWUzJF/I/u9Txy4jEA6xudWPmbYOTWai7a+2Fu5x0VFE59TEtPs9fGMVFH1x7uDyuy
afhHFoMKi+8Caztbcbv0vGmHfZgIK59boHf90TAcG+Hl+J/IKzooOgb0AqCwB5bZP/P6kKmRZzea
jzzKuOfnJgYpHPlclybMmH29nofXuQPiiIfPGqQ3B9Gd3s3Mj2fXEaINs1eJvS3ttu2LXLkKyclC
FFNzZ6mCJZEcbEzbipI9qpzSSy5v6eN5DcLAJMbe8eCpcZsqj1uNo0C4qF6twEsDUv/VvJXgChYp
uIr+x1bbkmsnpGfwI7AWaCadjBF6cTHwqii3hL0dKhmhQobTf9mjojFSIsp5jL/+wVd5De/qUsUg
xvChcFU/lH2xbC99Bxn/ko23Q5s9tih3TK4pleJ9isj4puAcYIHdX4f+0damQA6mB1CrlVOLt3DA
7RIgJmisp6LQ+aGEmk5YuYXSSazkjOlgwDYimHB/pAnxN6z9rOC+dIDq0GH7Zyx4e0ok1zX8KAM7
mhMf/je/na+m4vZuPRzrKpl+FbONAWFqB4+uFCRMk/v/yvlZ8iv4RpM641f+EozuJU2JRd3Yekb6
BUmBA4Le8IZmBn5LV4hd56WE4MMBO0VcVhj17CW0csKXzG0+ayk6kQa1Rm8ZSPX62luk8gx/gvzn
rJD8sbNMpuf1HBdzWrmfKONJVvafSESqWEWYcJ3H07JdXDfLpMdCedDIs0OCiZbYjCOFXj3DwSGR
IRJS8jgljpPB8+XKMiaDjUIl+zB5Ilr7indPY1W311lb6lrRsJAPpI4bowIYzuyNmU/v+w0CoCjm
Mur03GwJkj1J1AZ5UWkHvwZncPs/zXsKptvffZXtlmKGoBjhoJ+DwGDVeTnVVnqy5ujCnOSVV3Ph
JhyLx20b41XuvOJS7B3vVEqoXbJBnHiExTLGB5bBl9PX4G+B3z5/mMywEKUI4WCdc6+VzNCLHxX7
rERgePXRcJa5IMMfm6YLKB7RGIJaOA+nfa58CLH18nIELz4qE65TDlKXSEWRokNoj8SvvYDkogHG
KEZJnzG7WPkZB5UxSNFyurzGKuS41MbYzBh0y0pYoL4bDt5wk4kNBadQ01PMTc0zkbYFP6eHePkx
RSgRuqOc+nFgzkPUM3cLAvMQCzVmryMx+5hTYJhMx/UYZJV5A8PiyZXneMdR5WFNm0u6d1m9bx3p
SU3UQ5v/H41Fp2xJFJO01uO4ctubWNWTI2hoVuanQX9NWq5gD8WztPT/WTWv5aHGdzXsI3Y1FGxK
KmbTs4XREFQ0+TBSraZ72lpcyigHrYOJyXpbfUxwu5x5cDoQVBhvfHvZUB1bHkfkoDLBTdiDH8Jo
2Ntne/N2xBuYOhRBdpN3dcKBHQTFIwXFllboD+4tUVRf5HdeSZ44tPZW2ieYL9PzUpimgUnFDAaj
YQy8SKrgH3s8aIbkiB3KIktLOtP4XYUAAYAh3BGpXAvVn1MGEBIDWlNq/cC48xACqahQKRlULENY
SoLDsp3gm+Khr1GBK9s90WcBrQfCjO8CLgjmP4z8gNxWHM+oqBATteVZ+9cMAP1u3b7MOF1epzzh
PPD1aBCXEvu5nnv/rdQgI71BW+otEPDxvADKGReS0qNwqAAekh7CGbR+jdFDxX/sCOjl6JDDRCpn
/mOs+Fv7ehkMa3O0wDYpBtm6XDEmiXrc4KkIOjDq2OZXcZgaq64/kuxwI0H8/j80siJ0qN6ZOO2o
jRRgYgNDdagTp2XT5cBfA5Ui8C+8veDYqnu80O8vbOh22vkDxqSAjlatrv4EPjhWufJGDSVTi8vJ
ET3xgr8n37Ve+/TIddCZSdo27W90ZNJKYKbXqIyLs1vBq/h68735oluDnRST8DeBa37b7eUp/ivp
b4iVufuNOojICaRpzTFbF6UYDf4oGFt6lpLgpevn7OnhKgIFfAU9EfT2pT/xkSQzo5VRqYC4aT9j
mKv9kD09CiywqZ8okJjU2ZcbFygJQTQoJ1h9DE3CnPcIzJAXMoPHTRoVBgxzbapZZ8GdiGS1YAHn
IYGGruK1BNJbXx1ykC6loxr9IBSbqyOr0cywbMkDtma4oerjFqkcLqA0RMYOQmBu7lZRkJJ3bh19
n+KLv3MdPTXLckUapUP70IT83nObqntiWXnbJThSejW9bYyMx1ksCAEQZ23ma+dvZkbxghk7PW/7
mLorFx8deC9rfbfsy8Dk5fHWXxO/g+8PCb0x1jc9oy5+Eoy4sXlRZo5yC8ZWOYmS6wjiKyaNMIQI
byzVTc33b3GaUbXO9PDqFcG7uryR7q6vWO6qShuH6QfUjfijkRhvN4rImFzamA6YpC9C2IKsJ6LD
Lapn/WiM9OKHKn/tjbcQ3SiP5bxDq9MXDxbSDvLU9YgUGywmQ8Jjwul8f4wTD63aMD3faJD7AQjD
ZmivJ+28BUQ4DSpsBpIuxWzUIYfJB81NeRJwgldmDMpwftl3woUT9VAjN+cMtLi8dDOLb4EmGf0u
+jh2LF/vJ49MtCOYBfupHDqzy39u93tbIKl+J7cDD2mGW3ZecWNRvCA5Foa7fw//MgRcE79DWAWS
Bc4qOnTJ7hYpsk+muL/TvI4TeuDWvOPHIVm8Sizk3A6oXDZPArmWa6tytlBZZ678kddynykTixX6
aKyjoFaS6mB3MY7vUloeMVGUC8n85kzeAdmbxgorSkvxBp3Rozd/oW7SrXSIrAJY0YGT3RdZtKoz
Q3a1se0Cl2ln1rDe1IdboeX78/6lgBWeeZYaIAzJMjPNCzU9XbmXR/713x1D2d5iNxGdznXzsSkv
fwmnirue/KAJNdJpJKHFo+7iYwzN5kgtuYzbodJiHvkswSX1O8royliBlYXpP6rCTQkf4i5r3HDI
Ebd6ZX/GR26VzYzEnt/4o7343AtPHqAiWnK53iJh7bcG+Psawpg2qJ9vC7u4rdKWmeHDpRFCrV2+
cntpJ1v4fWvrMoJ9yV/GgKBhN8ykA6JTV1sZ4s9LA8jzcmgY+0kLIsGSsZE6KUNLu7SOFfJ2sWSs
SNro/gq01PB/Y7FZ+4oaFlBeOTvNPZIXvFeD0MiQQVr4R42TH3e0SrTCQU/WiV85EhwKoaaeg63p
yieWFAYgKWQNzSB8VQ9j2oXWb0rBBhfWfaN1+m1kfOmWBdlph822h3CNGhE5vhwHPrBYVwWnajDZ
dt0r+6Zmu4KajIGyq+9QcTiwHrEyUrb2kiBO3kAbQ+PZ8ieOhaN6pi7Y3+hB4WNPbMPb46xcWDUG
jYRypArniN8sGJBMCY+3p2hNre7vCmqtwiH5MAa+XBLLlS0pvcZriBmjkRqGv+GRUTq0j0svfsZe
nc3jhHwOyqq4Pt0Zi0WEJih30EXo+8Tw6YOQmkZy0XcYFlRGxAvgpzgj8IWPJvwNinuzR4YQRQIX
SXxj4d0qD0+mHgwOa2fH/hlSktt58i70N1AqcPXuA5DsZ4Dzc4GJXByX+8qsWRaoBw0sJOVg7S/4
OjEc6DLWUGRNmdb1oD/5ciieDOLvCYH8Qd2FXBeJMZ5z+OuzUXzrXge2gg3F0AYBwT4BhCsYy7PK
Lz6UT2DQd7IYUUGOp8O8HQmXjzux6CMtwUUhaH5WZ9wAPZMNL1hL8gxIwJozo5vQrSmTZu//0VWI
T7zpyIK9slkILywsdsyqtTSQmKfiKv+GchKkw+j0R/5zqTEa5hbh7TCbmbTrT6aJah0WAlGNKetV
boK2oGHwe9u+c9/JPBNdletoi3h5tWpj+Jm6+N8kgWg++6IdvveJ/DbfepBR14Y8ANyBtSrElu3e
6BOQuZJN6Z6Tys6GfH2zJLrsHBGOZ2OQQOT/MEPpbsHI0wYEodsUWOHwiElKYr9KtqukY0HRNIvi
gx/fHT1WOYF7azaAn5JZWCHXwm09bET6EaUgNss9mV/DSwIOuf579gW08qdGFH9mZZom5Y0nSNTN
t1EqKP3tY8W7ngDHScUQ5nscrd7QYfXlHP/OSwXZWfmIWewwXjRzJL8yUo4B8zpCwW3xwUetQyF3
whZnMWEqewNacZszPv69hjmls13oIcH6CCqC4TQxYHWuv4B/oF7TmnbdFm6pHZ1hD1Xn8Cn6BI0t
2myfeLiEgx6f2xM+yx/btuM5F7bIXblzSYu+u+kBd3RiPoL31TQS05bmf57J+j9J6kdff60a86mP
evND6t4bAzNwWHPqF3qzIYc8nxUCz+zocFvMKDKnjYCIMI82rBGnIQlSt+h1s/YE6nI3H4LydRnD
IU4II6a3DLQKMAsf4YTelUmNMGV+YZ2uwbR7Y9YGiP1VMBq+BrKQsGwX4Wapn1gm40caC31+bGeu
r2SNO1gC0FOyRQ3k6AN9dlpje8eGTGDvf8vNeJT9kLUPpUMe2/EOaND/CaBCEn0bOtjCdjssqPXI
n4+dbqnuRhv/c6zTtzXKMo8gFMMxd2wwfICABot7o5Ln0txsiM61/69ESoAc7JHHlWyoZe2RZYEW
f9XcqyX44xjZUwPAMgaPyBa/fN8VGHd2nXUzy99exzjYciceAaA+Z2kv2VK4jRVqopBluarS93fh
pbRQ9ugVohXIIWHb1so5J/zZ8/c5u/oqqymAUlru87mvMY+nbhjfVkzrfvbuhFGUH2DuV5h7zHpO
+VwxZw9Fbu57m03Gr6yed9zo0xKyGu6GXKTdhyPvFbfZ6rQlvUc4RnFlvOlQlgtqYNqLV5vsEC8K
8Bh6TQAFLWXgs8vixYTrvQJzU9s07N9m5XVp1XGSBneAtyTof4pitkeJ8ycmpHAj3ZNDj4BtQ1ib
2Z+29fJAQgyPQTx9LXKyX46s+wSfBX/mCe8nGpYl/kUJfscnfqX4gHeEWsxOYlVpMo1kiF42Mva/
LUASiiyP78NUpSSFROPAjLtdH+9BD0pQnUGeKEErjWcm8wXMm3/Y0she6UFGg0Hpf76PUVdMg44c
zQZxjM0TW9k/0cWY021eBSJpxLEORWz3khZf1K5HTlyB6yl2vNd1gMBGTSQNZgIC6e4+kcLX0kjm
ZtH4ljnWcQhSKX2DkK/SkTQv3Jm8kj+R9I2987WZdi91OEVcVY5YoVh74KnrEAPknnN/Tv4SD6oC
HDok544HgjsQjcNXfR2H8iFGb68EpC3qIWlDzlIaGmCnoqwrYDqNATPzmTfcKUCFsi7p023E5QFR
s8VLLvEXetQilIMkrJC2eSejc/mnRCDXS/M2WwvUjLPJ+OHQkNx/7XQe0w9m+icprasApNIrF56U
H7fFcpufQOMMtor7HYmrdQTpF8IVYq782tlh6GVHq/kf9RhC4Eep+oILDVlw5FYJYZgAEJSd1UFa
EVTdA8907hTAQsRjNheWSTm2JWH2VjmnbonrnXZWrk4+KW+tFHRu51T894HgPs3eTNxnBHZasyE2
P0XQQxpE8pv+GgIvp8ap+C9xWYjQKQnMW6G9XuGpWmYGDVaana3+Gc7NX6BSRTMzasHD9h4Vlxo1
i4BsTa3GSwMpU9H62PTtLGCjd+a+82EOXejjTwridSpMnLA0iCx0i+VoE4OFVz8VSO7wvgIiwxyY
ZY6XCJdp/RqetClAppRy/CAPEM9bLzaxWtEUP/mudx3j5+3Z/Wqk2qV7PwG21hOhN+azbYRqBWoP
rujpt0h4AShCDtouVDOdOcp/3+mjYNncKhyKecTQEcq7j2AEhs84L8OZz9JeNVrF7GZqQvz6lVQ1
dMsEV5KY00Ur4lWXR1Oc9Z/hyz5Luf7R7+A/kn6hmayxaRDJZ1lxphw/Mi8aWjETg6P3a5oNit7r
ftyy9dUpDxx4ySy46zojJ8Igv8U/b1AVUcFyhSPZRMlNQgNukhT+DJ6xOh3q8sU0fOmWRcB1w7OY
AtbyZ/sGrVasC8OR00IzZjR8XcvI0XikiC5u3ziLnfIhR5oRDUpo6c5VzwBhbLgQVSpPdEk+Vt/u
wY42iFAzK7C6Tz0+9ETp6n903xCazHjrkgsOItSwfZJEJVgrrXyedq8lw3CVqjAy7Nrq151GZcL2
I8fusFqa/FckSX8AOUoyHvOhKzVJzBPkK/MnT0dNKkqS6xx4T/R6VBCYEtOk1pjng2+c+WHJsrtP
5H4T9iF84PLmkpT/tgmTFA0WkPzF98E77MxXK/gcnn/0Fsudq/1gfFfpHnWoMvcc8vGPyJurJb8N
IPaWweKrV0GNDCat/U4foxkIueNvtMEYPWu24QxEDQaawTc+6d+QTBRyS+Xn4qjYoggfbWMqSg6j
dwnrr3nWeKTT36LEB4jJ44UXHaoAH1sH6ClB9JhG7sZdOMXwhMaAgFDSdUmkx/67+eiXYFwsdi5u
ei1dr9Of/Z/Kgy9OBqZhLoaj87wIJiXEWDwEiHBerdyjzw0FNKN0GtQgCF5u91dCzh4Jvhg640VL
SMXAmGbFf2ajt8TL+Cs7t43xUpiF4MVkWyA1ngnbW4KdJRdrifmFt7PL0HdEjuW+bdef82Iy20QT
ky74cv8P5JEAw+She5RMzg0MJgVntPM3sGVXXvU5l4zuroWlextxv2p2mm45NninJXx4G1HsZoLX
ZKLdGrvtVLbmiZF0mziBpumsCjFtjyM0LEPltlRWOhihmJt2rA7+O5j3k5dgay6y1mm7F7P99sXU
eY4Jehinmotb/cy49SPFfYsFHdCP4VvrtENJhxaeZV3abESO6+I1CuPKEGim4i/W/sMTnxxs7L3D
z/FFmVbFz1fSBhwcrus8m8ApSvFKzQOxrN+A1ZVxUpcDbIL6zd5+h6Wp7CbaOl0EeCU9XSpQzsaU
rAG2bOWaAQlQO1X9p43ZC0Rdu9BETsK/5jpauDv73NK95AclCVbdot6N8ddtSI8/NcUkrPKS9xp9
nE4tA0I7AfmlOlIrq9WsB7Wt5ZiglkLhFsoHWl1HUUVSckrL2pHDOpqEplFWXK2/VGqoTHC2ndq6
76PvasDRcJrTg8xfT4/BvXsHH1YWl796CEdy1//rtcISGqn8aEZ9gmz5/Kl5VzPLlfv2OxxH/HOV
WagVRiL3ciDVEh4eK6acll8D1Cmap2Zvl1bnWRZHHfim7HRLZ65qV2CoaBkBc5btFTci50pB+rLC
SyD4+H+zxlY0KrzvO9WwFkBYu6QOwrh6Hd8hTvFPnJOA4on+STwQnYQ1YYwH+CRXqtYNGTIcUGMr
WkZ1q26pXDVllwIvaUiv0xJll0vGJloQ8Vz4NA3jJoHCk511ukhXorMoatLTsnVUGCqRZiolaG2X
5KiAgMcD+QBUVDYLJ3uX8X/Dop4/SzCb64rPkHor4iB07fdnFhexApyTlZ8yVFStakYscksRk78w
F4oxm5HE0WESUzrp4y+Z0UwyV/AUHoybHeFNOo4nTvTKyKJ4ebVBCND9TMjfXZHXPTzaCTvfMsRG
wJb8aefxL4JpQw3arScl0f0LVtYOAhNTAdGschy/u0f+jlKGDdGhK9RBaC966kqchrQGOpTKPg7l
BVoL57wg0lZV8G3MaiSGIXSqd8Nt+O7EpoClpBNbUsL4xCw8UK16aEDFursVxJmwQOmvwPnegtqS
vAkXO5OOzUkl5T/rRGWho8ubZnJZiwjl2DZhR3WEhGySbE1DuClSh8S4H5+osfgGVSsoKio/ZVz/
07c5q+6NI1vk/Zs/l+qQpPGEJqah0nf1+6gIs2WfiRqtyrAUhCyGjYMXzMbaN6lJmSEONB/VN56F
mlK1i3AEp45bPeNYTI4Rrl0juc17UiJsIR/vhS1IFSSUNqzJ7DOly9ukcEXESPgD+IuVzYqBgNca
HReSH0TXVYnKKPjUj94EOKMKNtk5mx0ZOr3HlJrvVrWZL7lYOBCtQDnQ9cel/OWv8gEglTEhkPK5
w97n/A4TVEeMBJoVCO5LtrKNxmDCZEZNWFxXal1RGxxBIA1cI4HZB6NFUw6YTSaH9CftgslZYuMX
i1YLssDo2msTYwmhTZ22OJqSn6RXz6LsykmjX7QtWWeV9GzqwB2DeRxjZ1FYFl5SJ9NSpjDel1SE
QAfLNvi9g+JmaZ98w9gD/Ws/Vhh2yz3DJFrFHeHHyUmP3Bob8ktcQKQ4i2USOwCZ0nxIdv9DhmXo
2KtTsuHOZC43sePthhuJ0kgb0IBeDF6mAcWvKRE6LChKB2dIEmscCxkwM7k1cz0E+TO66KsYfP0l
+hmmg1f0OCxefZYeJDKC2RY0EiN6Co9cUPydrE1xJjx+qIUsBg2EJa9WmRno1HBqUAV68zKvWD08
5bcINPFINw3Zzwm4FJpDF0FQSaVmtDRdCHeiR9XS2mqkf6JwQja+y4EUSTnvjjTQ/bsiL0nZM234
dNHN/vFef3wZYeUzFL4s+sUB0cbuYymdYxoQfLSTpKtmNmjq+T2Emz+BnSMOYNHvfKafjZlHFJ7Z
jiOKkXvyaAZbRNh0xJyQX6/B5pOPQG+kVTASD/NF7oJZTz/Un09MTQxqitLVHYY9Ti0+UZ9KVvgz
zJat8tXWLf/2JNBK/GzCC9ERl1tNU9ajmDRaER/9OvKNEgfld0YlCwQcwnzNn5p+2sn1q+8Si5k4
IGbfdk5uiSFU5eHtvkCxo7PJLlxF9f75MM6p+SI0CzZzArZ4uMg+H5oX+UMLZyc/HbSvd9wFkh1v
3yFnI4QceUbcSXeEoWx8f5A2JRyjT9hgBMKZk5/BYRq5MgmG+4Np3469JZtKKNvCgq+wqBfGUrbj
OMenpOdp0syiY0tvg1Ee299spqPvGbY1xrwbXigRTl09PCcgR6Cc+xWgEzuWTIhWwRJt2LBhpyNa
R+zoMxr0X4xijnYfjY+EeZR5htegmaQieU6Qd2STCekwhW3dy2Zo+PT4vPWXhcJAwQI5oJ3k+HXJ
46hvRGgZoXag5SffENQW9TO+2+fl8HdkCM787jpKqYCZmRaafL8T5ZccQrCqtUA/W9tGrokLzAED
7FRCEfMWXMp/xxc80lNX/1Im+scJg/nkriAW3N+073mCJZllHECp1fKVeYDyJddEOr1m4j/fTYq0
2HZnEXAjJUyS6V4QXaoYMGhGinykoyj7vZcGg8beg1P3OOPqUrNLmVVzh5ZomxPO06SKYtVU3Ey6
NfiIFUgZdJacQLO3kAnI6ku5v0DYOtapVHrWIjgT8muClklymuXGdX/s9qRVpcO8NYoT+HcaucSF
P0nRL4Rd7Y1OyezQdydm78sFcUaZYgCPJ45KYgZk65BIgBGfUI6TZPyz7kOULvaKbjE8G8cFolxu
z0wQ+f3ovT2TPTWSQWEaDTZ44EgNlzr7mn5Z1dnQY6XtVhpckxl6eIsEz/pxIjQt+XKEfvG1g8sk
1RtXMa2/QZyIkHsQdjHmSi2eNmJSTuiktoCeeqKxgL3JtrdoebrcXOzTwyJcWRqDf7Z5Za8RjEzX
Oc9tDTIvevZEBA7QcZrFTJaBdzi7S5kWNAyl2eAzXy2DaGdsu9dghMbnnnr/iWq8kpAjBZ5ItJOW
7aO+P6AB8aeEPEaLbYCuo6kNB9KkVV9vrOn2hGvyvw2D8rWxJ8TymCzWZ9gNfivqUPTlfdYILQ4w
rtdr99zzU+gIbcEMJypiMyWgQSLm/5BGzEa/EqazeTkanq6tjpgm3o7KIBGfyLx9ChuivJDDXF/Z
uP6HM6CJb1YsrPRKscIBlW54lp1qNX5bTLGylOR0clec9D4RQC82FjxspthLgRKdf/DAGZ4yfZH1
LYXuUbIlrqjlTcQ302eH2Od/VnDlBRcGnAPX45CXpEmVt6++N3HTzhQF0Br80jlcdcaA6+0uJaq5
KiTWhD0/pLCaSvLuR+LRwEAYhcqFXBJUyakV0ZV+BELd9MHOj34uXOj31DpuUUgsnFlyKgzfFW3O
oclUX73URJcCBVq8vfYdwz2WLmCKUHzIP04nb75BNQvVfIMWG/FDHYjCTXUmIcL8tt2oEdROTYoM
wVW6+krot/mCVQJ+UoCZBUE0u3Av3UtGXcbhLU8sAwvAmWGUMQxlEdyKc1lBCEJMvsAqbIKXfa2P
90fIoT0bxNxkf92L+cjcXN4HFk0FVhK/9YFlWrktSR994XGtIkcWrcRkxkFS2/J0iXoqelAti8DM
2lKJ1xSjZRjE+3FJT5hYL1n1ii8xe32pvl74utVxmq1i+aKSr8JIaOgYRn0U8ntRUvyX+pH3fGCM
yMafLTAAbO8HB3pp/83daLrTf1D8803l/hwz+cze7l6QV9Nnxq8cD9hggCKWEoxGT0OxTjSNTkt/
gD6jlDHfgFrS1hZmb61Uc2F9TqcfynYTHwENz6aGZQGXgFd4IHW48zQYoY4W1SQpCcQQNdc/Vkl8
SvVa5SHZh+2xXLpaXmDPNQnUsNdmIMg/h1a/+SW+Hvoc3iR56HvZvmBYeLhyGB5B3fq46Oi+HEKS
hotMofhA7zldHcNqR0sKgL8MGGa183Nc4zjb+dSP4AucYzhEhVXpPuKeHne9DcL71+4zup5wc+VI
UXb5vVOOZLOiEuRzuYVyKT7ExqfxQUgK08x9/FCm50wRPdZ4Tedo5/3F3EgwwX/PJqflCm5CHjRd
G69HDAY2w4Ao3AZOkagFKHwiNl86fPFYYwbWACxV+c7T2nVxkIO0zMZBvsfJAX1EJfNmdjYW8ylv
2AhgaOLZhBQLuzsNf9qZJWAWq6YoTHv0sYY0dKMiMOCx756URB7wf34nvKAC80ttcWAec+7Agu1p
yyB6p7Y/r9u4CKLOoVMHhDD0UwktrQUuN8NdmGHvhXmxmRUPtEO3O+VCE89L/9wB05ZVo0KvNeGM
1gRUQsWh3qI+w00bJJpzU7faZrm+TMZ3jMBFOAmxXyOBrWoodwMCWqABwDKyH1Q/1qtDH7qZmwln
FUvfKCEvsyLtUzZRbQzXxXarfPyFbon9XP8zjsDw7raAMWRZ5kmVR7Vmwy9IxKZGLEayMH2p8da5
1Knm/JwCnFKtwLYc6CgkkDqeL+pQyMNcOOV/1XWsfjUhUW3N7bZFzU59HGSaUeNxmeRwCylm5WJH
wCrZSm8htsKZ02tmeA1UWbHJsGrrR9BQNrfH+YSq5+O8/40q/zm60EkN9mEKQtVo96cBgt1UFIqp
9hutN7YX1EBkZRQh/HYCls+bxRGj8oPentJX9Dfi5cKJkbAxzg68Qv42ywpQkTLk6HdGb3leZglv
XsO3gNkQdLw61h5ZKzObTJOBDUCq6NBTYWiWR4Lp3xVEJODY2hR90o60Ww6hSK2qZquXctyHvkxa
MILtMTYNKDO8utAyojRvdWJX9RoIbax1o5bvbpqM2tgYTQp8G90d9sViJyYcscCJjtRQpfEaircz
PlASJqiEGfmN2evqWST+bD/qarq+QLKsYb2B5EVw1ML0S/s2YkmWPaTpj0dliPYmIGe8K+HTivDA
EBnZ36f4Ral9JiNfS+8WPWWfVAy+y1fA4IxWMtE1h4DZozuhUImIucCM29C5CE27X0gNDGZEcGd9
VRKszlDzymB4DfzyWPnEyjWhu76jMxEFBG5mwU72ex5jxxkQ4EyWrT3FQPmq3IiMJAPJzLY/M40/
ngiruMth69kET5eHILxw80kzG3a4fxgzJtPE9lt7b3q5VtewvRicfWNW8W9MnNR08Zl8YIvoWLSb
NWVE2CosR94390gV9v8DxjTDKPaTb4k4ztvxhdIyo1AIUdY1H+99uwccxcqy67wMqyzD0R4wptg6
uGeapmIOFt950niiDJ5a3hrSOD/++dnpADsZU1jK0ZffJpHZb2QiF78BJmKEqTTmEDM84qbL1LFA
d/tkR0/Dj7tVnjrePca37kTKpDe3FQ9NKr279phb+LRSNvJVcvN7wZcscJesONIJzQ3fRwmsAwfE
h1BACKnLivXjAahTTgO0UqldExdtZIKDkz/9r0FW5hdwPHPDO2rkjjpHuHkav7Bxv92xLytuAvv+
K2baqRWKWYAPTAQ2KTV3V3M2PTEhokjkf2m7kLplSMjoHxkDiKfi8J5+JyfrSCIBet+OYCv/8mYq
osw3BNkNwsO4E6e7M99AUaUPGSc7XwYHruWgv8eAsRCXXioPwzzLbQnJR0FVBoa2u4LLYtyvJ1n8
mD5h/PFKnMV9HxtjpkZl3qHKDgTVccBde2HyuRDwIKVHf2nFDmFfrPi6xHt9rCtUki2P8W/NWZkS
j0yuyIVbTtNlD4+J3tS4raBtnU4T+2FZhiaCR51CWHoD+ofmBwbFB8wL3MK0TG7uCvlWam4n1JLy
bS7DIv+dE+0/ugJ1GRN7erUwj15XWiJMAaTl2Mkr5zkVs+cNZALnd4s954HLdo/HQkwhNksxbeb+
pl2cwZn1EqgOXqfwt7iTrnQSgvXP1FjLvzshbFv9KyaXqcKfO/d436OLPkTrZOD0zVbA94nMoyD8
E9aErFIMjzoyuXIt/kw1aEG+J/2bJG5oj1xtoIzRfoisgTMDIMn04sCm02Dg5qBmG4PWkNQI83Hc
z83v0J1E+tmMEkwYvlhpE+66ADxZAP28LJ3kYqFiThZZkh+CtWlk4F90hoHPElbJDZ1DNGN52sZg
R+akGV9IIi65vlTzEeCdk15Uby4UYVjDCbjtJcBcxm4vhXtSg5mHKlWR1BhWZyyRGFV0iyD+Sixm
5ONzR0EUkr7CTC4RRmRggXzVQppwcamX395VM5+wGlhjrLhTc2M7I4CB1x8nsb8zlOy6GogVIAYj
Abfh49zPeZzU48iB1OwkwwNkaJaP0GpNaE5/POTblkdwCy1ES3EREITPfGghs3Lvj29RrKei7G8Y
NkgrK0GnikPTkUV/Pu7id8SvYZkGRZ7MPjeQbFDl3yVnJN257VWucXczBkuG3gNhy2Y7QZRGCyw7
VD+g5sBySBcSGVgHfSYDS8a0ADvo24gHMrLdcSJhH63+I0KKIHVRuymWQbHoSEWp30qtbAHSzIlp
8lcoFoj5QzzQGMUm5dhIwyX+3sllZoo9yXUQVnERMF+YYz50Y882u3/NXs+UmNfixiPKZeG6HaO/
vQ9EtUcAlFhtPmcekpV9ehTd1xOWHjP+RyelAW3HvSVtQQMVUsV429Ldq0cEvtyGfh7NghffFpTj
ijg8uXJxkX/hO7ad67t9sFeKhoLP/IIVSCnklXEoZ7Rt4b31g2Plgf4vXwNTJoAkhxYI376Wa9g1
G6fHu9CeRo3VCvNEg/+5oXlbuIolLPpTwCR7rJb2YXLzAFm5ngLZoZ399lEWZe+VvhIjCnNqqpcn
elcrS7EAVpm105FNvQ/v65Nnk0SNPRnATSueNpoxoS4reyr5cpRzxzKWS3P//B5oXQWqlosEuDhW
02B9Ui+aDLPcbwTc8Sl2+S37CPZ28NFAiBZRiZhayp3qT5bnyBUvZxrgewVwfZZQXFtCB13gre+O
nv1AFBgbwLl2zwN6gkYs8rO/RgZuV0CFCQrkf/TJrXFXn8S4PL91sShpxnRBSR8UXzLh1MCdNgF8
0iJA7lUm9Uhid7Y7FLCbbbJnCHYwKJvVtkYpu88o+HhVMvsjmjUo4igIuiII4Ucjl7SR+UvP5DP+
RdSrwx5OAeTrMRMaofD9+rSM2ZHIEm6gPm0sBb9EZsUinf8OHqkMW4Vw8mN0EuBjO91WRvmwNX0S
5oJV/qZiOoHjJyhRu/iqnOTvG8Vu20SVkzjLmQ+JkMrpOf3zf5fsVcIjm1QxkMCrOi51IG0q1LAV
veOp1VYhRqI5N9TE553z6NMjh46s0FJyCvo4l20Q4fdIChlW44StivzkXQ+b1DtHs5izyntdNBTQ
TkwHwcs1O05G2tsIntSTuKZcDJvM2Vu4m/K0iuwpUmxNODJtcCQKP2mZLQ6Nzkjiwv1XPeIomL4H
CsTaf9IrugCf0PrglIsH3SC75HgM6wi8pCnsU0OvltLAxJXIJfhkTV4Iin9qcEmY3K+LFzwRLJ9u
CPOrdt0RyJpyvK9cfdhi5Hmot0KPW+JudpcJ/mRUyhk6wXElj8c5bb1CiKAFoRs6WBWx0UTckJGh
bqjlUI8bEroXUdno4MnYcKY5MoHJ7DIxUJ3NZEhU0SPOW0qDl55s+GzlYuRMgjtw1cG2JS+OFUph
pbZOAqyft1Ek2ZOHJNGe6v2czTVysDnmF61d2jwlRHJ6nCYccyD1gwnjJHWdkvr/qdPQb7OCrUnr
E/JyqlUSsvwaZqSJ9R8/5eFuSZwBE7uwJ1Yzs/0cRNYN5hDIaKRKELeHMJULXSC1/cr/DIrv9/R+
yEaBIfCeD+5VGLy3+CjRcABRr7sd3Y3VC10rMkpGMVSR3u21Nc2rvy0lP1uVANJlkpI4CTXzM2CM
hZhgEF1hAeuVSA7QawoU18Wn7YcZvBtxAk2x4UPlneXsW0u/fl4EUoIZc5vKjDug2/2m1lYk1Nsg
NQMvbRRoxTC4nR0DktEEBKkKWMHp8RUVF6jYhheaBxGegNldANp34HkHAfmnOUnwtcXg2lMIvAy7
jzzyqRpjxX6CR+vfh4qSQNUlubmIXOBxoYbekUk8uPlSpqTuEQxJNuooOn9vR/TThP/pzeDHGeap
WLAIpquFpJ4hEYPrdwyLS3UCd+h+Io84ru40Vp/YlYmaflKbyHE/G/qFhSZVJ0UaE44thUpS/eCc
Ml5ibcnuFNbY8Wy8cEOYg7dmKj5exNc/TvwezImEb7whKQOBPh0lQCn+N3Omedt7HgMKf9urbPCp
PABeq7zC6x0DtPNTSuGDkPq3owGBRjbloqIRgEtRsvp13qeOvWuqQdwvSDFShR9mAuNBaQCXpMFj
tpckE/0jHxREBMwWu9A28Eec8N5nzLyTcoB4M7SHCTfobZAe75tSsmBROeeIpxY5MQ+1uDdOlRl7
gr4LNx6PH6uv3dWdyeD1nDr7Dglmsz/HR+Aareee1PtwaUYWIf76uPBCODdPPMc8G2bCd1tATwio
SWNJ42CCWhVl2I1hM7X+KBP5Md5k4pcoc1ubKgdMYGXdCDiJlFAFlPTEa/AqKa8iC4d6WRzuTrl/
F61RDdizj64Jr1IheFHDhunN8hXfsVKEXI1CVZQYcx+iCPaCkRu8y5nEZgjr90St2C2oS645Duwi
SzVnaCLNMstXYt+pAnYdTNv7lABKO27jst2Dfup+6t6kAcZatpYJu/ibN5gSmO66RUrgwatKw6Je
XAGN4PlO0HbdDBfKCdudO2chrC/pHUMiA1ROSIP+dybAgUlzNH3WYSAC9xGPUhjWKe2qrZWmT4rC
8a9UJ5DNQmXLDyVUCs1b+PGlrZNziL7IoA9wwdKjha9pWJiPJVBJ65Zx9NXAjIcUTpAS/euF0v+g
cHKnIrycFuphIBlatToew8oU8HVkRx55BDKskDwkivjEC6vEv75fLg104ge8jvGEBJ8MKdl+uwaK
1wcicY/SIhHiN1b3XIbRn2mPTdrhYOef3iD3hF8qLA3PA6TrhuajHsQOM0fMZe5cJgEuRo17Pfc+
/0Lc28gfi4DGaothX2FzWi98D1C2oD6uE5p4l7k4162n0IJc/GriTHdT9uPseXr8v90qVGa/fuwr
OFswE9OADT48/aHX9AnPdlh84QOPseozqD/B9gCC/Cztho/zZawHW/nUprQSlRLs7jKbG2Stc+4f
+SmD/TW+yLI3EBfqvWG6l/7XNmRlvxaSBYWavadFZcQnkBn6NjteEUchbfsdBbsJcOqFfoGJ4V1Q
cywJKK7EXUVDouk8dX1354U0eYDMdjycqRNrCeHUG+IKAjs5j/RG+RcVvXCgLY/4pUHy4gFHSKFe
6gK3EHmUWISNfSif6mdWKEEBBAD1U5sBH8xhgsh5ZHXJFV+3C9FLsTQiHmUzTZtC8QnILHq+38vg
8xNaBpZb78IzANaMCYyyrbN4wjWRoL7LFgynm3aMW55sm2Pic+/UyqHSlyN3JEOoQqrws2R6PeTP
v7G4an4JzmrrXgG2dyCBfxW9PRCmdpRh7U496hCvkhaY3IFWq3kxlgtwRMTu+TDrYZZ0kQp+VMKA
58uUFrFMXrjtDP0pmm7g31JOpEAr+KiT9T/qs9crDt7wVfvAiCEUgi2I/Ny3momanDEHju5M0zjI
eydAKf08ED5wSkGJYXkKnNMwNafQMqXwthks4U55gv1PIQKZ80XCHEkUXjOgU29ZE/nZXtZYchCe
amknd3Ai8XdfnEUHOCAI/UHtFTk0mVjQJ7NPGGh9gJ+3zeJ6ELC6+Asb0yOYn5F4nHjKUONexBwp
A9ernA45eS+8OLmyz++mZaotn2HsS6c+KPnyK/LFZmN/37ZUpg7VjmI9qD7OcLeXvewoX5tBVaaQ
/Ctj9fj3iZCzoja+2/yIaNaoJlHjy/oo4CyWY1ykcCCVq3Wj7Gm7HH0afp2nxpz3kwjhzb9NNMws
9520ehSEOiskEk83UAl8DeO2jHEVAQNW7ATz5GXIywdoY8l0peJWv8evZdEa6YmJr0gX5+s1sklA
q/Z+RqX+i0mfEVwVATcrLo7QU3qMUjZiAvuE6D3EdsCP7OXvJikXBtP+tdN8BI1nqN0yfaFxVPD5
0gT6tsaZct1iygBImYNuCRyvV0qH9WkgoBnp3x5hAeqODiyoK6cdb/SXeKiU/rL8NgHB8yxdI3cv
kEflz8xrVXaE9xuqbX1p2Vzr3ma6xtYiv7gGesVGyGcahL0RdtvLC5BnnKi9FY4sexPDbP3X6jrj
xkQj05JJQvaaw77/3Ev9tdbVv5FpRp888pW/ndhIM8iGGxyeW6kUYgd73RZOHhbGEOaZ4105M5/h
f1wlbGohD6gd9NLtydcjV1VyatDY2AJYvmPeGTXsiSgrI3q6PZbN6sa7wgUaWdrg/rYAbqJSo9aV
0unjookmVsYGW+M87644zEEI3BIAuO0llkRWiHxGu+8xLnL26Ce1Py0n4pM4Zx41PlA+9YtDm+Qr
ARN8Irpng+VWLcN9xJuEqyJeIC6rm33+25QkU5IbM2NAwxgiRKYqOYgHltNSQ6REv6j0nxwaNWFF
EEDHvvuuJiTbKlAj0IfkFu7Gr7smccgbFggibG3HgGydW7y8vtTVumqgL0iXDxSXJD1EaLEWNB+C
3BkCmoiKZOVaEYLMxkqvUxpLuPw5OLlRESdjyc3RZeGMmmxgcAgPVTGnbYuWd4IzQ1WW/uYxhynk
QVXBDTNwaw7hcuP6xPGia9v8g/U7TEMKaVmfba+kG9U3OlYpM9zCfEORjqwXPPKLmW8yxDi8ZlKo
nRURXDlx5CkWrRUyLIUf7Wgt0/k0mF4Pyr6jIovWuZf3xfRT9ui2URudXQynaPngrHfGufoxQY02
H863g7UzoI9C2NfuDh6980apVISPfbwi5DLB8EJswxOGuB0c+cIdFRIJVYX1WXf1t1JiQJ9+cpZA
IwAlz+OZkM4Ez95BqPDvO/vZfSfFIL8UZ/lSTKEVrS8do5/4U7jrQ298BC8DwKCTUfoAgsP88gUm
G1lKD6GbDtz/J1DKEr2WV1Tc9FQPVMqwI8hd7oTbt/L0wbsic1rQ2Jf6IEgM/cZ9N6nt/vNQVQO6
QQ3F7FiUSxN+gfMseGZ0x1EaymZoRQ9KQGoUeBGrYqVY/90f7XYsRLFkoqi0Pofp/STSUX0Ln60N
ouX5WZma4Ra+5/Mcccxjb6UYbY73JSvwwnBsbN5wkba4WnR+Pn+mw8hcFgPUDSd4+eEfrOw3shU0
GbS+0k6RW88RjIKfDb+1gfa5kt4KzTpGR6uokEuD/czqdiiK04BhciKfRk49+09eXKfQBM8DzypG
VQQVZAz6YAblcGleC7VkRXj8W69O1EfQMyvOWGvys15w0qJ1dlWXjyydKE7a4fAIfJO/TF1xYXPM
1zxI8egbeo7VvZeAcI/xlsOcf3EK43+Wi1FfiNHvpkrmQ+0Apqfbd0KIPyncocMkY6t5PqM/DOBf
N8mErWq8b0k2kpVBy8xNthEXPQKODHSj6ssDBF7wsnMckQfXU7BANFBAfjo0i/GwLEUPhKYWvWaU
GGFh+HhiSZDwEKSb+4H3T5ODMostq2QaudcJmCE5Mt0TQNSuAWcQnyMGR9ng2ZZr4HrKfwZNQyOM
thzAbcOWgvKngik2wpRcebxhwib0XFoHq4XuW8Xfo3W4TsLAZixDBdMhi43ifQA04Qy4/6P8zBAL
ZUEYmRBqUlhgvUxe/v9xU3Z40z6UeEx40w6o/stRCaPszBmc+ZvX99gy0o3koXS/yipE6iSWe0i/
HXPbrPCQnES3jmTtXHCHhC4j0gYBsVq9Vc0vSa1+IW2Pf31ZzqQNuQ/KrFH2UZCMiQEhqqDqjnJ+
k/fxXknp+TeV2//IEP63FxizKKYu5OiV9dM7PiBMc6PD6EC/QG4qrEgzAHPJY0EedYTC8+jiyJXT
u9pMxJzWwfjgN+KY2LqhIsYHgN3AutU1kobJFKNQRd8Ztfi+iuA+rZmCUQn0x2u5NHSaeHxOyUMt
5Qz2xFDXG3I9E0CKOKt7NyGO61R5pW+xVjmxDlqjOvT1JLcZEMl5asuZngAdMmqBeDqAvyRY4To4
UbBKMixDKl3B/pOSkONUswJwYnqFnYeJDgK2cNDSkiyutcPARMcZSHUMTIDYdfgExtd8HJBpXLxI
vMwmXKRgeBOKul871p2zzcvFhUjySCVjWB2TbUl0Cv2hghQpVhfCS3ICLL2eRj6aTJEc7yRe8o2Y
b3ykxChDyq3cjzS/0gLHZ6CTNA6sbTQkinuZ9CWRJMIU1hyfqtkGfrxng3B6tYmj3Js/2qOUnwze
up+6Q4WJyBkGOr5fZ1GHgmNnx7o3C4pZ6+TNGXbctpSV6wHWx7kzJya/zubwzZPEcuulXJuUkhzk
99MMsq2Iqk5trJrN7/6wDaxuEzgGo/SlfP7KP+xSHI6L268cxc5uHB1rDo3Fg2fXdq/NiO1n36xD
e8eXETTKPqf+QR8cCD7veOgEwrQWCCS5jGpl+HFH36+/P5np/ZySMjAt+cAy60h7QJ4TxEZAdE3b
cPAqc8KCxveLruup4W6xeDF0EaKURUJbkeXWdsV2b3dvjIC568zPb46RO85vpF/fcx90z4FOZy3T
1UmipLEUSxH30RUYE9mEVhpScglE9t43inFd2NrAzqLkIhiRi1P6W6dc/3iB61ulrAcDP+VEHTKd
imaTIr+6ne1dHdTrrcADobornA/0n35TccXlTNGnQH2TeBg0NuOeQzD9j3NAZnGDCRmOyDbzUAA4
OBISRwMHG5RqkUKXV348Ho0sbcoYBvW9O95oMZhJIG/OL/UQu6P02UXYwXsZS79PRzRrBho9pMfI
4VeZ8zy703cbTXAXXRG71BAoNuePtKOL+Q8bCkZ0jFfQv+LmwgqejyuSDFa9UZmSb1HuE3OvUBDG
8UAQ5mMRlx3Ga2OEPl6DAH9ksWEQBoRfF1U1Gh+2/WNd0dnBk86aHfrMMFx4VLsmh1DpLdsjtriO
ERklG5xFBMzoZFgBioNsPQMg6osvcn/T/9sxjlb+NtGoxVkdDVaeF4LfHV+1o4FkKQZj+/gQ+GXD
2Oj441+DNEHb47k/vXPzd//4E8Y9JjtvriptQjiubdOzVLLpauONsCAeqmh85KtKiKQZSS32vguH
HuH5h1xagV63Rzntwe8xbB1Opa3KPpwnTAtQN01sOdhNQQKYW0DvYdfv+Y5pzTdS9RZBcOxRFeQP
qhYbZ4+5YF1S6zK/vYYKPXXbXA4KXlEpbEguTJ+btJDEwehBDlOnfu7TGkBIa52jOO8hzMOqwdPQ
Z3Pv/eiQIf5vyZ4KB0MeRfCd+xNkpXtp9Z0uGNXe1J340Qk9GNHV/5cdjcQezWiounTRjORnft9P
+weMBunxJjtMAsnU+pP83v+9r4CoG9UllehV93eE86nxHWq6bNQcdpX3uCsfCXScMQ8lB27T28uP
wV8vXJwzz1Ro2Z2rAcWOUdyvwvlPAlVDHfjb+eUdLgvyH3/UsuEXUGVHzoPky/hwym7/9+VAb5Je
MKoX+zxo0xDkk2sfvtNysCE/xmeiqM6j9xcrZNQ9vspo3LCRUwtirBytLoD74yS5dfdieBnQAAVb
UdaIraC9iq4OV65U/Md8Oel4Q/I+qhuDXAIAGjnXAOhLkYl3BC8aI2/2CrBwIg49GhbQvGILmyJu
qSGqqjkpdL/6yX8/Szvqs3l8gfqa/39ACyFLex7Kba1M6RndWRNBKxPmeNdTe6IRdX+Ie8uxP0QY
bvr8Bc60N+w7Kj3xNFd2x9qnMQZnQO/VPJRo03kS/ZXEOWzSiTtLsB0HR7sLvcaa9ZncsEFB8PiK
ZxO5St4x/VGmIr2AdcS9Ob/5jgv1aY9O0ramf7Gd+jmpdATPLk3Nxn5+g9lTwKCKrVWNMgVLv/+J
O+mLk/UKAxhg7D1Etz7SPAZDXeZLsJUpoezdfQKRG6tFzJu6QSlh39C9H2oH82yy5hZVnBxlV0my
Au6XDskbNSCVHqC+/mNk3Xza283DASakcJG9oDpNozb+0mvKLQ1Ghb9mawd9H9SIB/H24UnwWpcw
5KwUhAP0MySpRh3xEXAvmluntsww8v03V197M9qNEzlZkh4bVdgWMa+Zo7iyI/+pmQdZhjDsnk2/
hwFfYteSVpOnnno+cDUGZCcu5hDueHJZ6+FoMpXxKKSn+PlbVJ14/eGwml4YLHM5D4dGmNz32Vs6
YyxfFJwEUO4BMOWkAGZc4mFu7enmVr3NJhfSBFvCv7MELZqCsySpxMXfbMF9IsXfvXFQrNkwD62S
9NC1hvhd2K/8s/NtfecF01TEdQ5QfNoBMJ9lCnJRisOzFhIdhO/8mx/bCj2f6ZbvqbWCcy/lxPd8
0sVOHJJioUGbJBu14qkbgcxRqIkohr13a3ynkCJVkLb34z0ehzuka6K0ibYNKsOALU0Oz7S2unBo
smTM8x+qxIiC9grFP+bNfD1mpU1/4EGIjsIQgMmYdIGx7jJBzeXFtzeBoFgmv/6D6S2W6v3nhvpA
T5KkElbuXrjMxTp2T7DVa2ep6ACDOrX54gmnCWPXz0y5Kqn8ZVywrLqa/njDNG6BmR/sUgGDhh9l
fv9eVRGezVMUwvHB/607B4sUbeUw0G5DIBAtQrn/gcKUpHRW9f4mpBhRxSHTBqpU9pozgjfrFtU0
gH7+oHW1FOuRAWDl/cxh1JlGd1WpICUp41vGa3xQjzaIBTAJOTItu+0UaSND33dvPLt3XGpTeHnO
wRgWy0/vWQMR+3rDGxB/kZvGDf6IrUttdTAg9nnxmgZ3DVMUZ2jct7K+ZWoi1nuD/fG8RbjH2yq1
+9Apa7aYQZfTHzUHfFpXvHrjAX+dquo5w7KDXZzAzQYt+CYyoF9/05XvgBLGGTOSVm+YmtorW9Fr
mGW0lvrS4Wmc4TR/TOSMywZT9mdhkzcnhpnMEOhbNk0YhM95IpmvmuX2mM+jsNMTdHo1uBIN45Ov
0GOm9bT349uigjUFw4/WnM7NeOgTc5D6pJv7E8x2PEvfHt1irp8hiXDcoS4jikL9YAh/2kJVy4NX
T2IaQ9Eeot4zBYQn2HQtySR1IITAejyUT4/toXbSiyBVmjZLVay0VtDK4UcY3bQbvTCfVMiWVjBm
EGOEhi5/UvLPIX9Zi0PKYuk2baRQLQpZqK36Ct8GuIpNRtDMyOZqzzHrsbLwxACO0j19kNZHbNxa
4Ldl0R1r8M/XX56CyQQ/8H1VPS/IpLaOnuuSW/DOodnNJvYXu62Dt0Dd5g6jevhEMEHiRAEKj+ZE
5Y5otqjL0+VMpeYqSr/OlaPaTPIIa8gFNXjiqfANN15dttXnxpB48ncaWxIXxKHjLbtZ9wwFVQWj
mF8OyJ8sciyNOz04rbKG8BDiU01MP7FNuxABGqo5Jd1X+mIzVaR1o84idmvnenWWOCy1RtGFumFt
/mg+dIHcucTUPebpqKBdcnKMyMArQIaCoIm03U+ySQzJ2gY5z2ZVH8fnwiL3Mro4Ba88LcaMaWbE
jfFfpwUdY55PU+5UABdlWItAD54R2FzFuFZCG+koJA/fiS0EIwVwt0epbqVtLF0NJyE1lGKkDDW2
CwsXHKtnN/SJegE5Xawz5yxA1vtn8zvfWJiIrAbgg8i85vOOyThLsdzbGhLbS6NwyJkCNyC19Tb2
iS1NwuwHeTj4z7vaokqYppRC50kwXDjdzDuEKp6Pk/8TjlPpkYummzLnD77PdWaaUxGi44sXRlK0
K3V8ASYew8Xvgt5vFa14enHbx5QGazh7M+qS9GIa3kO6bL9fU9vahUDM5XljtM3oR/dkDqlg5iKo
Zz24n5C5mT4H26busVE9djwWlKVikNK6J10g/uhzHxsYW7kxLXXEXKMT0k0FMPo1ZhcUa63vHPHq
nBdToArG9cU2K1G8RpBL24Tkj3gSSeaqKf49NG9t5AEGIq8e0AUbA4VI6wg35d9GdW1cQhlI07Mm
sS6sz/s5VQMbDaN/K+PzeCZpBzHF0x8kUZmQnFXDgGljyypeVEkZVSUYwXxXko0c6ZB5RGqKaFpi
Iag8Q5Vg+sn0aQFy3dUKjAf9EjrLSikX82yZSb5YJtopjSH+WlmzSqzdsUJ8p1coXo2JjDdwKEu9
FQTYcM6AR0zJWrcEqNNIslyKnJAyr7/6dvyaAedrsG8mQ2/BlI9rGL7H+ujk2z8IrIr8sWilimLg
4eBwhMcMrexBrzdMKRV77F5NuLWDyw8gQA3KGsXG0PtXrLuh9CwCL/LTa1/V55LyZ4L3HN9GmzXC
yPN5QsdWI/E1GGEWrqGXCNe3mkV3CCChdRrX2JLkGh9suX9cBYeumq8xmHgNutcteIr49VEosT7J
OP4/2YK6n4gmPGTEmYUe2h5me8qB19+zMT2JXDrBU3lNgI4MYSTdipNzX/OduyPXNmIBEluAoiy7
ZPV9U1Bnn50kzIRWSIhCs4sk1+xGMYlW0lHZKbc2TxwChoExE0XkaPIeDReTmmR1m7PibVtBjSsV
jJ5PQLn0OKY06OeAidYdPHQm26eQsiiSAihu98xZlcUSBMWFg749n8X4H/VZsjd6zd3BT3ZS4l+L
r7gELwiiKVYr5x3PkbZ0sUsa7aIXz2U1AkQ2FxTyBGJAgjEfiStWs9bvLVpSTKZYSA5S0iNintkE
VOh+HljM63Wk9EKW+61+pNFJfFaiTR0lzrHhhus/mYgNlo8CCymDd69XtExkiEwUf79By+mDgoHA
tzAQaWepsDGqOZ3DF399JA9GvLDbEhp5GpcBDcqjLgzFWSPr7c7k7mNOKuVJU+OLknbdvQHDPoL5
rZx+PZi+sUlazIjlHxQELiXxDXgjNMwyCpjHflfgDXEPI6UqLofW1dRWPSPwLUY3yhFK44vPZsjB
56/yenED0iSDBdOcL8wOOMyWiTXE9bog59W4obQqoVKdoSTuJmVCjOKFQu5qfv+odBlQhvZYN/al
+WW2jG4SYMtlJGz26jxR2jqc16zm1swTMW5tILrGawkbXdMEJdDnCAjtt+sY3Q2UJ2XRHIx9Q1up
JMWAAoFUozYu/32862rRE/EyOV+GNZHdeYs1lnCtiJyZv7eUf1tz0fihj75m64VX7g95vSpizL6O
gANvYsAy9dg8BFSVgiQ8jiTQ2GL8YIZTxLv6xAn+Rdr+tB3H5x8mg1MVLRpaOUlS0uPev39DAz8i
KByVdr+nridmHkaDyHGt50CXuG220xdR7cyKtueWNLH5jWohTYrvM83Hz4hgAAiWftgGNP959Fbh
vHu0qXvCIfVwzJAT0Lla0QhvxCpZ1n00tnaA2LiQqF6R+jKxVDtnw9qMiLQXFtdEr25iWn5UkRkR
/VCP3We6QEbqMhDUXPNXhnCpR0eh+5XZW7yHWbwJbV1kk5yU0I2qUPvgBXr+wlw12X/gwuYojLSu
cQIEIOgT9+qi6ZWzHw0y44pG1p+/SkJnkFBAhGJqvQW6/0kYE36/X5TqPNuxsWaTmqcL30AXStke
c1Vx7wJJLdhHFDknqUPN38zEwz6u8Z8GEhx3QKiZQFc+Qq1bRfkojkAxYw4NoK3kSMSoV5ME/IQZ
zC17HRihsSc1GG1dgLBU1Oajnhak/Qp+RLJdm5x1P10Zjg3RS+3KfBdyC54v/wIeCLmGVV7MLm+f
UjSKTJwkS/rzj8XiYBU4aDL9A4mLxXfQ2CE8WbTdazyoLjg87ZU6ptmcoppj2lgp/63XDGHfl+nl
UBs+0a3VzX4/UH5KRIqFeQE4MyBIq3M0x1GmRaXtoPfnMUsgO7JD10RVdCwwEd+yqwSTz02pho2s
BFuunhq56mdc4zqyLtfQovdK8AUL8ZbXXt6//F8+TbWF44Xm/zVLoG0stf4ko5vPbbgcr+Zwi2bs
pHwXiXaeG/iWIKFcerroWTY2sup+S+8NqnwfLOwjZ4HdJe013rMjJdXAf5vJVw/iJbRMCjKmyAOs
3kRvx3GwLu/Zwt9TpHwsR6l8H3bpBtPSYfBZFSWhbECqgyLNGBkguwMfW89F9CG1OJRXnp3YUsp4
VdmHFGxt5XiJvesJdy9isdT5tL/mYxEHpsdcdUYnqU4c9uwZBk+8LuA4bR7SXE0iT0A9yHGr2x/U
TaKzqOaWeuUuszcUbg+mxMgq7Nei7Bx4FDFBcdspalPIPmtSllccmNIJBev7JztRgEnaXxqJix1n
zSLEhnl6hs5yoPlRGAH1OO+przCeUyrkKNtsBCq88emHQECuliIsmkf8H5677vgCJJCkZlvkUkl4
4hLR1oOz2ZGzg+IsClX+hutjrabaAoTOWpOq3G25ohnC4UyZ6nJd7EuDYOPv8xfYLhAf7a570MOu
JJnpzFTO5qSNqNKYCpR50SeKkW5IDK8tjUU6JRLXJ+ZMhk5MDN8cwtygEdC9/CT4ke8dadZ99LUk
C3PAivvhkOLrLVVPA1LmBLVBdbI1BMR3d/+mMU4tn4iDF8ACuQu+tRDNcRasmehPsIvAu4xyePmN
aAHEY5/EryCDyxNHwc+Ut+xhjTp92j7jPJFKe2w9qd4EjJ9KBzHf0mpap65YX4l1hoQUqNXUCm4u
w531iRHnjibjJrdLV/aIPGNxsrGKNm0yQjw+m5okSeNKGokYp6j7s7ODk8x19zNKFCb8TOb/p+fN
+djUNd0ZyRzUQM1xNl1wbMZF+0hxSRw6/iqNKq7+l+luM9B8mxPdo9KH/SYKomnoFTaAEqZnqn4g
bZJtbsycobSQCKv9ae4efb1qzkZzsDGdsmW19RQsLrPaRoDeLPudWPBAnER1V4LP3BblJqtiR162
/prB0MOZc40n0jhwJT2iSHlPm8oFFRqIpu0mhUbcMShYFCwx74L+bw8AxINJQ4+774JNelP/49h5
Y5mj4/eYAmNgY7YDofIJodfJpLnyFoXME87xaAvkCvBMW3PqWpvRlRAytBOAcAbhUtlvYPH3GmE3
5nYR9wD3V3o8Vm5dY94vwyuWIIg36kLr5LYO8poqqF6i5+R2zAtytLDU82H1JgvQkrvTG2llGGBu
NZQT+pVYLR92whcMBF2zosEY3ypgffu0Fd5onxtQEgM9Btq8J+sK/zVc7p3oHrrYzYI0vqhmThJ/
EYlxtmTgoOArA9Op4NFAdV1ZaLrggEQrRGK3DrBnxJdjTFFg2b99oMaJSD171fi5T4pKl6DvhNyE
0n2lBGkLkq1JAjoQCYgRq7n+ejHFfRgsByUKIZ+7D2IhGtfV7aShqeckDfJwKfLEfJlEM6qtqxW/
n+Fh/fLkpr1QWSYydsyufsblrX8KqUEUKDUU+hYyz0YtPXmAfGlDMK6psXS+siGG5K8GZC0K41E9
EM5ORNNJcJkvQ5PR4lQ525QcglfBj5aBay07gJe2lZusOF9IHTGufVcvtgu+N+mm18y2qCKplozw
I0rUr3SToGdBK0KND/Tsujhx6b2+KAT2QQ6PzYHHRXI+tJe6K7F/qnp0CESnzIHQLdw8UelpY2w4
JxkGyayOrTz2u9OJ5fpZVVa7460iMoUp2gI+wz9EpbkFmaFo4t+DVGylmZd9gYgJ5yyfmnLt5DV3
G/vvTu9Z644pg/gDHbdk57Xot5Nc48zJX7+9IsnzPkp4kLS/B8qfNCcOY9lcav9qdYAmKbETpyBY
7Ws2kh7MxJ92BY7a7H3sCAcQkHLTgGiqdiXFCeNTqwgbuvbVk9NATtve0QTFr3YK1sOcBeJg0L/D
VHbgXlbBi8Z9fVURDLC43FBkeJDC4Yks07HR/5CGU7h14zoTgQTLrHPO2HTHbpWURIlDxJFUMoIR
23+4pqIljuVbI3KfAeaJYRTbBEUWsGvIs1IqqlJbIdx4yQZk8PJPJd4dmrrIVJBh6UBOoT0yCc3R
sk5iB0NL2G1ISKRc2y2bR4eP13YGKD4zhwSVJge047OmA9ZPbpKUTBpTaAoiFHe9XEwcoka+qtZF
whpoKbSH2nq3MMluPSliYQpsVUMwFi5uqoUgl49CKCQi+5O+N5C2ayxGoTgNTX0rD/D0ItAiZYLK
v8aOoOU9OEEnukx3Za6LYS73ec8X32gcEKirQ4g39eS/EL5EwcAGQnY5li263axKfnxURqQ9QlWK
Zi1AI0waVVy07ZIDFlbLOUcTWeObihkjB3FkZmuKdjXQU20CdIR/STc+YbGAROzhQhERDwLJpsOl
lSVDW2JNHO90VsVr++pEC8PN8w01Zf3qCVcQ8F6u7dUb66o6sDf8oeHgZIhomNT5AZkViyQqnwYS
EqnpkhIl4Oe80/s8CN7fKX+5L6zm7XNGQeGx+l5gDkZe2b0Bqklak6GBdASwG5AfIlG0bq8Es4hs
U/LAo2AjvISayfKZvfw68FTX3FMg2phAAgHy559pT8R9hllELgl7kFoR0q+Yt/TlGEGeES68Qs7r
uIqFrXK4NKcElby8/FfOszOVzNAEk3EpV01G5lSfxAs9I7AnwJmNz+xPa6k5ylUo6QB7W1k+NeDb
xryUSY92WoNckw69Abj/F61oy2eRgqZAPcYpFTxCiCEMtVzvo9B7d3SkXitDYVnfDZ9LryvDbDVu
xRfwV7P9GYF7AZMUKJmgLdNbq4TOFu2aTyx+I9/IFAYujqzh0fXgsK1clyWYo9qixlZpBBZzXjQQ
h0ji8FkeeHs1EiWAeXNF8GQT2B8C68sAjhnhtBHdlJZ5GuRm/aGmef2h+N29r1g3j58EcEhnZ4gV
Djfl2HXTcKwLWgkpbehyxn58sF1FCOjznKRADWwpttrp5mn/3KCFXvSKOekk4HbAtaaT6v/g1yRs
DKEiZLHlumpGZ03+R/v7BIdE07zaH1HEJkjME0aVjYgE6DBS92qiyuh5pW7+ooISbhLEiGxaSCkR
jDyjwAEArblQyTXQI3FEuKRmwShdAHyZBt6OqFR1kpN/gJdp6Dau0hLahrWFoY7KKCZrn3ySYaa0
KAq+E4fNP6WwUcgVn8eYGwAvEMmkn/xZxOuJkk/1bCGbGzzKBNktPxZ/+oRFBjE5GxhZnS6OFxIB
XmiYW14PGcgFUb8+OXTxyEtVrYS/MiffDsYDIn5B4FVVh5IKfhlVNkBzz+sCeuHImtsH7icSVhgC
Kokqosv/Xa1GkG1c49pZekI/FoQseQa8sE2ZbG9ZYlfEijQja4s2HKdTUbzrFFFS+rZpn/PbB/S+
t0BETWzf7w+w34Twxm9tF+6qoRzMYPF3xhZ0J6xSc+F+wvJU2Xp851vgOsrX8/XMXShz75V3Bxro
OdPGbhHqYen5DhupPls+D9UVS1iecmM9ymjufz2fzH/M3JYi5jF3lznNVzdy3pCn1m/Y4pLoof1G
EtHaEVJRB7CZ1foRgvy6ubqKN1pWw+kDsN4oSd2AH6E1E/4/xebYnxgeMhj14bUvVZEUaxkLQ6nk
18WlLN0QXU6LIkQz0L1dUJTYyoJki8g78NunA1E+QblV17hnhBR2WxXClelGguDxYgfz6JGJ8TrE
wRjk8uNgFbk1gd9obZaj8DDM+JnvQLool0daf2KQUhg+ICA5jZsXEODUNE2zCPn42uMHt/MienEI
wzjhD+u2CCzIW9ggCSR9XqJVfK7bxpqvLVEfVtaW8QynxO1zFvzceF8aJCJwJMW8U8f3tfPgyiDj
41c6dKgWrxouCSUunT94fAaBEPyF7ysq4/Ga8tr86qNM27kgm944fWHXWQc7d7H09PZ22qCq4wcM
Owe4btLP8OCPkyHP/FZ0ML+XDldB3neQfxVAwcpettIx4UzQX2yq2NLUGRBGUehZuBlUMqlzFY6g
hgWnyBoBT1fLA8szGaGcoeZeib1KCphofSU/0QWIblrOOBmssIQCQsW/+1hgnFQf38XZqOrWQH9R
YjXKasSuhD9pIeA17qm+MzXK0n1q6Jz6qTT72F/QZOa+GXeo1EhGgNv0R6xfrFEHXHpDrizkwu9g
d39pNHz0rJFCwNybc8Rq86NKoAP87S8G7n4BS++7ASlQDZZgskhbmxE2qk7tFYgXg4rFXFkqn3py
b09heQFQyTVL51zRNAKIrXNr74dHnbF2CbKtEHtlFpzNPjqPcwA2vBGVMGHTRk36iu60t1Xc3luU
y8rf87CP9DaczNyvNR4plp+MEUJ+Dbycz/EygHuH6pXJ6FlVszaOtN6SQ1NEn85HUc/btxQ8g9Zj
iRrcea3x3DVfV55Zc5hwrP7VEMvk3j1VRac7ue7Uc1KRfikyd/6g6BOxGxJUC4EYjIYQ0weEJsOq
qb5YWWQO6sr0cQQaBY52nY1jEuuSD0Yba6As3GS1b9y+jWQvUqWGy16kF/+3TrNC/aorYJHZpUYC
O+O8+yo1u4laaKjrD4IyTHuV3l9dYqeHXIRM2cUtMt2TV053Lp6zV4Cpk+ivWeWbz5dafflI97Ar
hcihfTF7AOED5yhkpLqynMBdPLYRJPUn1Ccd8D3popilU6Nwmx0P189rqa7BiCLJbtcApF5ZEB0B
GU9vVakF+RhFjLYN/8dQlaTSGNTvtumNwbaHGLP5pn/OqZshaNjPvotyDkLvJc+ZlyF1nnizD4p2
4XZ+V9CXzt8BmNUL7pPsAofWE8Eik+0PoDnyhmXNNvTS9L+9STS187zNKQUG/ZiZLkqo1K5C0O53
BagvajLi2S4kNn35mzXaZbqENooMdeU2qSGtypXrdB3RRdFGdwpp358bK6gFQSLm08ErTSk41Ymh
iY4pR2NaIVBYDL2kWO/DKyeyqDqS+zCfMP7j0/MZBwvr2O4lsvAhzaFH+PgzPzggdHWAobGLvybe
jBXMSQQLcQ+9lziAq/PfJupiicFrH2YaxpxSaSITLJLLxc71h2ATLpFzb2zPtkPQAKd7/LRUuopa
+igVfaMNLOP9v4qU4NGbwWSJ/+YE1omTV3Lor3imoEqUBEVcLMBkUcr8wjTasmq2m8D2ctIWM+r/
gihct51MfE+HWXAzss4WtZe6LdWq5He4XmgRJq8L5utZOXMpGxb4QTdt5kzI1cPQIVHLpul4OfLZ
AWR1qCYft/0+YjSh/0QOxSdb5hiasAQNxqjOgHPXRgVYCxFAD+jLuorXV+LR9lxx+6b4P0C3zz6J
GUCA4FPECef3fEJaYvj0z/zGNNCcV1cPHw68GUFsb2ac8O/Hukg+sPDNktN6ZibZouf/Wwnhw5kd
9oK/UXxHcXsGvD5E5bFPvWAvQpFqJEEelAKHEa8mEvXC9Hi5DfwFu+UnDi7W3g9lro8o0pofp8nr
gZRF6tqVcZZaSvVorIX8KWta99gIdyQkRcG8m+Q8F5EP4D3e2udf8LO1u1wqKNA1Q16YwTpd/IDA
NRJzb2TDklJDzkB+g6azpEjtKx2Ffd5GxaWXd+PV4myp4kIzYBN2invLmAzj5lwZQzH5l8+AnZ5C
TiInb3rl8EEbLYCB1yJcjC6eHpE7lRuUjvwizDetDCPJeX5XDaLzAeiEZmzrrEypJNFue+YfTrtF
uZJV7jZYX6S8Mt/c0qc5hKQYqPuUkV4zTqbhGi0TtRwvV3rqK9B+7yuGH0Xo77XKcZNIC0Z0EOQu
/8LIDG8Wj34tg47LF8m2uTL3ps4+lPEWrUrOCVS1ZHD1hHwv51JJo4ND/2t/ZKKyzxjG1qRbu74+
0u3zvgH6WJdzGa0ASdAjYwDOBRuta+dfZSSBnRrmJBvYVBQo6Ahqe0Dh/+7Khb/xoP3oLLCyo7kn
YA9ns6G5VFzEhKgFGHRv3mxG4KN5LeYk0yp6QA8SgA/pBoRe/vusACc3HC6h5ykt+BX3dDL2VVTR
eL/Unca7hfcfnLmodq18HBuT+K8rB3agyt0CvjiouqVMbRcmGeECgUhfH1lbsZtA2urNYOaA8kG8
nSGt+7oDSKgLgnIzXiPp1ItLuCJtZsGThBWgYVMk+dViNSZkig2sUfcXVA3Vrq7pjtboa+p0/2tr
Bc4WWCUkQWEP731mlHHINIog6aMm1WJbqneU/iNuD4qj6rPjlmh+w0C57noYx9TLpkR8FgKZyLX3
NrpTlGN7AaZN3jLoX7iW4jkgK62tDxzFr7Vs+KaT03oyVYxBdxGXTpLurEf0Ur78t/Bl0JFZCDVU
eYhAvJctX71tdRFGA5MDVOn8Z7EuLcuwMmf4+BC4gi61ccVeOe9BNNNNIqETYvy3mUBILr1gLjPm
CmzpXUvxXRtJbaQ0kWNwXCKozLVtkqpTzwZNV8N5yUeUZqHWfpnkncvbjqvSplEb8rukdhHeRSv6
/LsucNV/LVbNAh5KvosUflVFGTbtM454JS2q7wJ7yzss9aAe2TkIbdyd6LcWvCBRYc2wORgxvE4w
GAaDx0NwK75eLMe7c0miuyBsj9cj8l6EEPBwqRFYmfBWPV/pEiBL3U+BZAj1OD9y4tjOU/KEBBhj
2K10oPfWaylFlnOEBKtdtYRIjLVqDp0ElpR8yNCLv9Lgki8S3Qx19gD1lPIkseEdna0Ko0OeFhf+
+aqzPXuxtr2zRgArF3QTUWTdZ77aPBRhFRKmzANVPnvnM3/lvs5Y1+QIXm3cJnM/dKqOM5GbNxFX
VjsiPcsgtIgZ4buznJO9r3DkbhoD9oyqJKSPxoptZ5nITYIk8mJF09h0tWlBo/enBpkBq4P1KDl/
mvuddUbAyWqtrR7kipPEEICoT/3s/mCpF3UGzLcTIHMWCI8j6P7lvSBjnfQfPDQsBy26OVljvEO1
plVnk4Xjp5fxkblsCSg2sYp79hNAKho2pDmveFeviIWI/8htVk2MViyIgHSSe6fF0h7T9r09ch1F
oSFDIxsMQzW/HT7J01mok6XTaig50kFwNENKHlbfuvAOeed6aylKpGps9UvgraoDM/cpDcM7bJUn
Wfjz0D8A8ej9osgqOxZqIuT3r8gZR4l0Jhl7r54VNZOnJ+78kWtsANo7lb/cSNXk6ylGV9+eKkB7
zLquY17ko6qMb1MvLbajcEUe0ILR7uMfHq6bFwIo9qkcFZ9d7PTgQ/FellGjCEUZdvvm7Ho8bNQG
VJib6jZSSBIgxbbLLzJjCIwaZRAFZ8Zo7QH43J5Dqk3Z3+ldH6fLu2/zghXArSF/9oZBewkT2Qtf
ep2tKLU5IcWTuv8mbRELNBwQb9Crhie2Z0ocsOGZOBaC2B4h/AwhiaKfIjltUlGfbZhmIt5Yznh0
8XHPTIKqyQ7nYtVDoVOZDOPJAYvjctfQ4L5mAGjzmrjIq5cEk1Rm063J+YhXDZmAx4vvqSOUDZjF
j/Hi2BgwRNj6mtwhJfuSeMneMVeWUJ+EQuahrNpiExVTGNMZYB49k4aycASQ5XhrOxgCE7sWSRnH
azqLY7f/lJIEGHN4ksyONPGjYC4hGLcOYQezhnleiPSzTYQYDIrrXPoOHd6NDDHkbZdqsmeTupzp
IB1dEil+AQYR7cBEAwHniA2G4/ilgkYgk21c/it7/kHXWw/Rm8nFbnAFxFcaWAFq8LjYaCHGCJ3a
ZFdxvMwkzi5zkZj1x8OkK71Gpu7uz0NhGsXU6+e4gzBP2DfqPrW24qrW744vCKIel+89RbCq41uO
BgQ+1E/8GtdD+qe0Wh06jr4DH8d6dv7KvcryG2ilzRKk7kMWYWpDCao6b8oAZpB+93R3sGFihQGE
wRV4EvME+c3p9YdoHFX/pr5at8iLM8xYTjKDF45+Fb6MeVCZyr4thsyMj8vIgEOR69RBMHIeyok2
RnNrRAFwfzSSgRuw9+LR2fiEBPULtvamVVfnAgt/zDbVpe2MYTqubx2Q8mw0VrvNiHkcaWwDsXS9
a97SzjlZMZteOnTv+UkFvVlGcQy7o8iyrIPcovDrGM+wn2Hb9FzAJ7huXpJms5ICcOz57kmyajis
aO2KmCDtfJLAtrf5edyFG206yJEtB6gc1Fv9Fe9P377Z6a1ISEd/qu6F3uMdVJx2i6f4tf90P6cX
AFa8wo+xLgfUZG/WuKeIwMnnf9Hwz4RwU5BhzJyEsQ+MizUWfApFoks2z2XY/cW+AxLwo2YVvSEe
UHexMQwQ18Z46F7VaHpBbhu24YqzaWRg/s+dYTPIFngNR5CjNbT5zcqOAylJjIB7DjtHFQl7oX5B
GYx3oNlrs6dS6qWeLFDiqHwTQCm5qdnDFETEIJXc+j/I2dUbWZvVAdpYo01y4yyCLiEY56ch/XEF
K+J0U47rEw3uL+FzWrvfaN1F70jjywYe/3pnNs0npz7UVQzyj6XzO02C/Bf5bWzxPBhCP5YoEbx7
s+5MebT2SvCsH3xE+cJ6T2P9NMjX4GSA7HPuxs3VzGUA3WNl4cBGcb98IHV3I0AX3fI/dNlIMgiU
zWM69jy3bY2NokMWNFNnL/c15eoybdXOkSyLtci6ggDbMHwRPo1mbd7AZCTFm/xtvw8BLyWIsrkM
nTXQEzCeDd30DLgA6vKRS5/fTP0lslgks44AV0KFboRF1b/c2KysskqP5ibKacQQYb85PA1L1gGC
kSAj6qMwFFQtcT9zP1HNqIkKPndR5XKX559rO1Ew1vX6nevdeMlBL10owFPT5N5Ei43DXYSJ6T3L
xRDq3D5zabhV0RXxbhkRNbVQZphpMSolVF2Y3M80LpB5cxYFuWxytPlsjy2iZiu23mE3WxrLgzht
RQsxJ8D0+zWKM4dJgI59exz4m1q1BDZxYWXBxFYVtFRftUNeEXzvU08TYDgUI1u17sIlDRFXA6JN
s5EC3h6KsXbSBG8oooxECTV0gaEHFlDNH88k8bZbNNDQKhiOIOXM5JhcaMHpTkudZ96Df2XXYjhd
0ARhnl9zlM0BMopqYTH7GiI56j5cEsOrq268BNKNHQ9rccPMYDVDwBOpSZ4ceyfQYvOaIVlA2Cqq
0rsc/QJDvDtx93l+YGK//Ir97Pm37dFmMBP+bwVCiZYNiGDqunrzBkh7cX23XcnZ/0i+R1xgHqx5
o5Smu2HhLRWCBsOVwfzVGF91Jwc7aoYI2S4wReAqOt5BHRtn0XwCMwnAsPQfvjG/ZB9TIWBNrt1N
XRIzGlKaXF9zBzcbIUd6Xb7RI9XtVQTGnIkv9AZTmxQuMm2MBP2ZyFDHKMzj2nFvsEhMmJOzpt9y
axi9RLYxLcgE8IJU3pdqipEXXjqQHeHg3uB2fjV56JSliMkO3GQSbysex2lqV3EwdJwJcuD1nMCA
bNipFEXoxYaELT5rSfbeQDESg0Wnq4kXlmg5lFyNUrCNJ/ry8CIkY38yVdPcYcHsoB0Cq4XJrpA2
8faWmcPCbk0JIMxAkgWsoPbauixFOMmUhD1q9ZLTaQhsYdSaq5V+DApNl3wMN7jJF7aUvlAMjyPb
7SqXdXERnLFR5cFGbFyjiHjruj/LCDXjPuSOJ+JrUEwO26dkc6sBE/YAbTscqW4be0HzcVnqGK90
LtfW++w4KII3UmttiqnDc4IAobY8x8ptU/iIOuo0fLuikDLpMZ5PIAQqEskBSq0DtNNHPc1sdvAG
ANw8rVd+uhou3W6PfzWr00IqBtQMrlgcxpy37qY7lWxL0nDItaP3/+2IrlibCxxgmqm9PiL89oxn
Czk2w0ipJy9bQBBCQRVhUA7zMgGpXzXVJkRdtcmt4rNMQyDGc+b1S1n5afiiSDG94A71E1IQTjki
l9qsj798VXMGn0FGqzpjNha2uXGbLZhH32Z9BAjJ7FiYjxIIWReZW8e5VUw+7ztky0L1m24v6+T1
1v3xIgkuo/KQFjj6XkJpmjMOO959/RRkz3QWjntisbzFztTVEhhBl/WzA+RuIS7RwBGMO57vGWrt
TmgrlWa07zPMKRsIFvb3F4TWfg1zSxmaS0ZdEqsSxyuMcr03/5GNv/j4WSH8hvZ10WQL0a/rXDKU
dz3Om7kTavreBVfWniv/CRU5MA4B3kP0Mhop0led3t9YVnkGvr75rlzeFk2KY5PSmt7Z3x7nN7KF
qAYZGt+F/H/lXFlDhL9FK/ARX+2vVSVc4oSYlUF/dK6HGT3qMxuNuoiJyD4LMvBep/xXB3AGmgje
tsJe5PinypXgKj9I2h/oO5p3QLVG0sRbnHEHvZq56KIg9ckfzHZrRKGDLdQSs86Lg6+CFpZUANpR
s2CTnIIVABUwGEKjZRHiGmAJEhPtQ2nMPsLUKSrFfSQnXHrXnqEeQg7gB3PbU77fAqMmLaEbJxVK
kQaQzvtGR7taxAfx00jAzUD13gkXlpY+xvuc1h/O3qpwji9VSEYhyiieqW9pXti28HEMqyFVFpqz
Ir9swT69IbblS6NlUixF72VvJ3WudMjxga3OHCWcgkzLoGHq4jFaayZWvDt4+QTLo/NOdkH2zd9M
kHT98vUAH6eEdifBihuKAGUmvdDCHCsNFLDArmokHFE0bOn2leRFYXXmg4JrJqR9m0q0tYojsOi+
4ECZSwniH3ugkg0YEuCOgP53NKQlUXKwpbH7ydLn2kq74u60QdZnqrcaEZz+KN1PwF2LU4hmhOyE
RGODz3T+YU7paEBkgzaAdK7a9mYxpQQrJ9+nGGXtLbZmO0wHoYsQC1sksoX9krEDd87GrlRE8p/A
vtEYkEJmKtAUUwPI1uMhcWBHIKFQ1KLBUptQDRrEDYER2/xaxcbwsgVpiCea/Qw+zgmQVuji8LY9
Pcf2ViW3Dy1t8g/UFzFSKLXm3k5+Fz+jPkXca1TIIumfxgasMTI8X81QgdcBqlrWaxP+PLeloFGS
FaG1PpY5R0MF3rYETj/D6p43rT6lzuZLhZrxlYAQR6nq7TpkPIY6NNnBst/uy6QNnAYm4mTai/hy
+VvjYe8c1n8yU99VKuyg1iY6NXK4iXPuQy5S/HsNG7n53ghHPVsQQMY0v0Ngs/eoE9iM3bmYDHcK
9RnkMM/yB6XPK6diqCt7r07DGYnSeA8zLtE6PTGNtQmYmFaCPSUfi/ctfJJbgEIb+Z+IoRdhBWPa
kKosMJWYI2DGNzSnC+jM1AkU1MifkNY0t3g6VqTjMd7QFIgX9uliHGIotVzVHatzqHaaGTrFi+D7
4b/huALpTP+tr01raeQLSD/6wxutcMVYRGYyuhoP3QsuCPIaotSFK5nOVWhK2CYug9Z/nQYrYtTp
IOJnM4sVQuTH1aIMNSBGKfsYdq7O94NVL1JEex0X3nIBd7jHhzm26oJj4ZqnnsR3rt0+m2njflwR
n0j7ORI/VSstAnuzIOKCctAzoPb7V0LTa6FJl+VGDsfBUyrKdgI8IS/uXESkRNUpnDJ/cVtmaWFp
gnwYgCa/IgJOM9kp71xPgKT7wEbrPmqV++3PgzHIpbo3i3r6VmGotEF74kqY0MOrJ9b3sFZeMyOR
2rD2pqA4NjFv9Bno56bXIyAGgH6FcKiveADOTdt8DT9/jwLFRkAYX1K9KTDLRC26SXuUgb/mNQBN
mNjMfbgJTPo7Va8tb1AgwIebIgNAOZXSkAdFHh5hg9Xsu31v5ywsSPBBNFaXRsZ+HNrDKQvtEF/1
gM9bn4BfC3ukBdtC2ssTvHQ0tc0FGuMBjS7/BdSzKq0L1wFotIQ6xOx65ovRzlQFCgzHRIpLlobj
fYC4lAJzFNqysx1Fq69r1xLbEGXsXk40Ri3O61iqf+ULApZdOfS8I/0n87SM2yoypjpE4D9conBQ
Hx5QZICBvns4l9Im/64wjlnY0DKO2xVoBtnSFvkM5BvC2baw7xP/nKJPpH6EnKq2/l+qVHlyU4WF
ALtIVXv4TtW3h70A40ISXOSVSRvXtHEU95hmpP21eKPWJo+j8WM6o3wqsHtcbFapQz9DLQAGjgPZ
FLe96ypQiYMiMK/WPVCBgkWX1g+aYMjv9PjG272Pe6enfRHWSb1QhQKKPstVpbZkdB6EfC07vtvk
NVidMIM7DVhgLU3D+/kUVEpvTBKQIgKsF5f2k3bczHBeg4FJsgEl0GL0plUgH3/07Sm17xDJRY8+
3G0lHow5VLi8xIgeRvOVaa0BXww4Jn4X68dxvywlIOP4HMowrNxqEH+peJkTfdTN7XpQunjZlzkH
mnvO56etv16SYpT35MiycCTlGdX0GdR61lnJ3QUL0Ef2/kX4DvPAC1hHxU3AXqnJmRZJuhjZDHxI
WoEPivg42SBFqa8NhEm1TaVVg6iz1UUAiiTbCHv1Qm7+4kuQb/5nvn+BLPi9S10my+xKihm2JR/R
IX2lszSgQ0KNra3fxpuslsDunzGTxGzeTC6WNg5fs2YhJS2wkFExziwgxGaBsuifov9T0H6e/F2g
3LtcQToKclVe55GyH+iC4ZxIwb+mvRK6Rkq9AN2uweFIUm0SJOpVLIO7yopQ7k3zM4X8IYbvQa9q
PP2hcaolwmOhEzKDagUDenrlrDE/kcTmzeeSaqBLCJwZZc0BfILl7Sc9nDvX1E0Z4PrFXFJkz1V7
dEf3OtQ8fySjy2TsD5ng04XPp8TCO1g6K2ajX4Es34zWPgl21/+NaJD6Tq+1DGfFn1eq3SKobNFv
wEtR2mIJCTVdggVJ6JPDPYzms1GyNar+qkIShsLZHCRJmlZaIzBqt5ZQVuYaONHRharct4NNrTyQ
B7r6+6u/vIRrtJ+W785buFXZpY0sNi2XED4uuxYDf0/TmcJQ4EJKcNQp5XIKLG107az5U/dhZwav
+praiRMqQKkJP2qpaut3+dHbD4iTLZ22qt01XdCDthPrppNXaFCP0uFUDCXLzPwP8PW1m9k2JP5u
PBb3nRrW1SGJZTDYI8DVp/ZtkpOfgoySEIonDA5ZYtFejHWZZDpbKLFy/B2LfdbIaKGESXYvX+E3
zE8okkGdwdNaU2gj2eTIrqmXXznA6Y3BQ5WzXYdyyPDkNkeZGiZP+2pCdFbx+l8iQyVKSmdrWjgC
9DuLb11H8/CYlIxMAX//ca/7f2FWj+JB6BEBd0jfY05DjNtn0lMiVD2d9iVZtHOZ3qPZdojTVQjB
vLNu5R5WiSeROKGVqwKR04eH7Wq/kDaLAlSGsTRlYsFDkSA/dVPJ35Mwh4WgrLoNEnfo9+Qz8Ef7
jtWNx/S/G3+sJftCeQvCh5YpSmvh1o8xe4k577eaokOodIcdJk5gJCu1qc0p/Esn3Y056yeUDDWo
MQEx5JZlbHc+OS4JWZ9Pl5P9+lDQ1QpaWPloNKSs7wJ+8BtCF3ellV73vF2UXMWZAExc8H9trCUU
cEyel0YWDi/nq76id9rZpacGpQr4CJil3NAaQQk4WnW2y/nuRCr1oZ+mTphzmjD/++cXxdYSSBX1
XNe1SYbKUv35UmE3ixP5aMTG8gTc/85zIsnyeJn1SdTK4Bk5Ym4xrFnXp8j4MlHfRclhhlRVqe2I
EYm2guV31CZV9d1K18H9ESAQJ49dtncZRlq3vidkqhp4zLouBEqj32BR0e31XlmVZlDPGdXTIkEY
E6ewrV/L8xuyiDnwlVwtAEdnwZoKC+tg0O84KBaK//iWJxh1X9mOn+uxG4cmJ62rnwudeJ3z5PWV
HDRldBdwzbT1eI57UQ9PH5Rw52WixqOFNrlD2ZNYkL7YSCX3OgOW2NjdH6goiQtQhWZlNH1pQhEk
4lv/uo5xdDbqypqvr6O5rToLv/0PWbenOOjypXGKS0D5d+YpUOas/b1TIAk/YS9ywBBUYoe9dQVw
VwyBMg3McXtmBQ3NlOflMjabQqwMZ4cjsEzqpS2vNWi5I3qdO0K3e/lZiqXPyU7SHu9wl6HsWWG+
8Dqe/iq6nbUarZkF4zOpKAU5yZcwoqsb7ouGn5fJ7taJ252mHxhiwHQsyRAMpxZFJc5LH82R0VsX
CND/0wi0ktThes+duvJfYdBOvnGftO8LcPbticOP/TLpneevBnbKhIcO904L2B2um5yZUznBZySv
AQMWOIeEIgKzdYiGNBNlQlGs52UEg5KRZg6Ep0daTqXMaSpHMJMLpv2LTNGW4s6J1xFVDhKrEtrS
vnxLDPLMYxN246QMgfzNeYtoDLqA+ItJQY18vyQk0SUkP4No6KlYwdsqb+DnqAU+Jhp+6PZs8cwh
C0fS1cjMFPRTUQF2agaIs0bNuOzZCkLucqIbQ5wliQmgStXHolkJ5fWRNS/6+GVrEZUIcr9tuoyI
QJlEpRP/puE00Q244UHLGm2fJ8mnonsJL+HNuDEeHFJbvlCqTHxw/mJu+BEeNRSEVjeX++Sf6Fz8
gm/gH8XkYAJYy1E8RziKMv5qTkchMmkRL+ccBMoc/Z5IdiMrR19/BJapseqwQpdyfiHBR2aigFaI
9psazhjEgTjh9wJ3NBmFHsCz6MO6rXuyin0Hmc1exCMe7mJ1LpeDrbVIxhcdxJw8QBjbUB/yHMP0
DOzczvOll4jjZEEYciCZdHL5W1JqqlZbEGnacFI5KopHdlKLjdztEM2KCZK3QERLdVoN/KKalW78
dEL7JUQpyCXXaYi2YzWk3O4QMmg3eWF4DCcxX50wfeQy8mGQBLZ+yE+f8TuodAktBBjkv51PYvbM
PWubMBbWZzwEtGohccG+ayNskQXHR5czxjTBRwUARixAeRE/LqMPzCgTFQ1BesUqeBNglaoG/8Rc
eHZbQBC0ifMPWdQ3/flt8O6u6aMXoMfAeQ+vxEft/75vV517mT8XTXAgQIQ+/3sM2hSebM89qalk
/jL6T+j5OIk+g1Ftb9W5AUmhgNtw5YQmqezQzV1zAjPA0cHjr9uTtLopoWgRvH0bnNyIRvzxG5ew
iUSw53dICC8vHPRdU6W6PWvp6M2R0tHuc0k7bTNZcmswZfX2/1puQkhEgWl1Uh0/cI8/GRyRfmOF
NerVqVanYZqZwF+36c7YPMwrqCoDKGLYY2CRGvNWlwthukufKy8vQT2E61oFP1OYS59iZUDUupFJ
de0WBKWm8T0DW/YY6dvURZ+vv3UsOb4edh07WasH542MrXETzkxmSKVwHkftIdCAf1I3HGAjgbLx
BZgyhnZoy1veHGOlsGz30gNtkUTIPvI+f+7hnizO37l2LzcuSbr5yG/epbJA0yKXlzGkyKwi5Hyw
7FegWxvP3G91drQlNr6FqnKwPoAl8HA4O4g3uAEfB00EdVMHWiVLgNolqRnxoHR5+UMJa7+uUWXE
8vqhj3l7fpCLvJI4dJkWw/MlIM/fgeE8zLT34VJd0MS33amp4AntVeJcLdq6+brv1wS75Lfqp/CV
x1KihsTBbN+n5X15BewtmEh50OlCA6F8LceUJlQyTzOoXcKoic9lD1X6C8c5e1e5oJQP2P/Te+2v
p1QtYfVMDcIaSzGgh4N7h9A2i5uzjP6r7qBgXr3o98wHWLGZfsCfj/VkZARBm2Tv+fCyGA+iubxr
lEQNjxLBMDhZ08lxEyxHBMtZM0XW/j0VSgdRdl/0k+WlaMFlDGB/AQ7i5o8knsYu4NS5GlTJvX1Y
cVaeAIrhDGmclzeD0m70Ub4PZ62x8fduIlJd72iUlZj+BeE2n6SeS/qufXvfW5KB4SBJQ1cIkALf
WG5r8gyAh4CJwGkuKriPadX5uxA+Qjf4BmokVuT47ViqyJ8rvAvmJwMRxDhxCeJg4+ULrCh3Nvit
n5L/hJVFwpzSercDlvt1JqouXC1HA+33W90tuBU40XrcpINEqy4q7tZqvTItju/iyAPEeEJgDBFH
buQwjC2BcENBDC+LVlQ3j0Z7DcEkbZPwcSuWXX28ZvEpkBcS7W+f8LFBXr3CffDT3q1NqcKKTlGY
SOYRrOCQ4jrtUC3hdqIzE3+xnszMwv9whP7GV8W8h/3ovWLYi65SeooTAoQSX3BiqjuBktyD3BvD
l6kt487iIheTIbWK6kDgH0SgFkzpRlKwLUxjZ5T42fIXcxxuf5UKh9RKg/uxXbDEVwwzUvPfgxBL
0MzOqFpKgr424GFmWgPsN2dWw9Ax2FyUvUHJXsSQAH5Pkud29lfcd9j1Vk/436tLDzANntzXkvMK
vss5YQJW2XxzsEZr7iM5mjYQ9sHqFlojoNFwxCVjXZaSjalSdu8vrdjfioUviShVchgTzB4F4Ik4
dsuRL+1QTJWkFc6qYEkpXAZbHNAy2a4FuM6tGJzcLMq5x/jQbTTlmwnYah4uWJCKi/CvTgWBNls8
qUfDGkxFxdxAdwGIWf0o5BjEeifDSJPCslShHSUlihccEcIlxylGgwEelsabAzRSmBpK7xoDB/Bo
e44F/hWSrfqMx8VWgZfZZw5cme9nc98U3O6/3Z66iubAdOEmUmxjG8Q8cABRULyu41I2TDfeuidK
KuIcjMaDynNX1s60LwjIMIASgZXdg319T0ca/UNa6FnHWfC4MC0WRKbAp2/Axf1woA33Vcf7f6rl
LC7jKkm3WjvJePU6tToGpB1W1Vxb3zFMHPlMTY18OJfnvQRej8M0bTaT4b1LOknWo26AxjGMrPX0
HSz/14L3eD7YuqO3gWfHvGuUoBzkCscmKEjL67d2rDS0k6hsuzUMlF9bYtLxfXRsbDo5Jp48Xy9J
v77oa/hn1pPMyuEgyTbs6QmQBLQyc7nlzaQrxsq+8QOgal7rZMAhRl+8R0TToGFGsCO+ZgqzKYHb
nwnVI0gYcXDPdyJEZUkS+DREfKchdL+NfdSQZ6dK3e8xV9lo3vmHW82+H+FkiC64ZEonBkeyyG8P
zuBZxl3oAucoIKrRURVVJyO27bipnarv1bgrAtwg0IKuuwQqfsnRrCS4ritQRc7RAm7YB3rDQogl
Cxa15ISIttUUV0CZwQDmXGgVkyobncKzRPX8osBZZ/RFIXwTYrFVy+onrCePo+uEUDiHbJmRBhAo
rirUdZL7rypbbOcsucR85lvEdmHFwi2JThOCmEVqK2lyXavimu17Mdab18hlZAig9Ql/GMWzYqo7
nCDcqCuJn4aB1SOGWZ9WYJtoGoKP3EJW8Vf6rlL7tfJV8bmiIpzr675BzKQNH5WHqOFwomAhgfSD
x0/7QBlZu0G0eOLN44M3M+FWg5xI8TH33rVNjAoLuOuEYT6ColyIW7gxUWwI8PfUpPlvJIk0Dsk+
6rojlaOIsRE3myDzivhBKsU7BgETkQuOe2rfO8PH2HRiVvu8VxpD1c1TdJEcqApfOeLsRhsGZHul
Uzm03Wdu2qf++m0Uc0FB/mu0UXsM3K/5Je+KrKeVMpzu0wybisiFcNxz+5ALDCOXCE+E6KKfVKzi
zjVSlEr6+k20Lzw360z17E69cUiOBKuwvZEWGr4E+hlqTQMftNfQXswDs4EHRsd1ei8TrHmiGzxi
FimKoAVj3xaZDydBavVIX6OdFxrKgSF9aNQXF/0Qqm/bJDOdERWF5xq9vsYdZofRZKG2h4Sip4rI
93QSPpe7nxNrgdIWhBOjzDFcyidutaXLKt3bWMYmcXar+J5qivuCihganOkfrV7/U75/zsQjkUJq
ulprqf6zAM/b5mK44VNem7z3S0iH/L4ueom+nwP3lOFblR6S9G3cSNfnFBbgW0xFB9AVxH3xPGJC
paTcsGNnfUKj/8JSh0Vji6xX1CN6xauXrfgVnsSfihfKoZhcfhWxiemmQHTKhFjjY6BYl5vxIYKy
1BETYkhlzthqzA6LgzKv0dJGYNRKJ9p7/bV4vHWVkg8IS7pZSsElZ87KaCGOKOxoRDvruCIiBxHa
qmeeCExrUOO7UqfWZ8hRXVCvG8ttMKPrFLIJN5/bCCbCBgJxOLEG+L/MqFvPGwslh8MCHax7KPTC
PR8lu5gGpcUoADEOOC5kF8JLFABYpJ9RkaaCCjPbcCoBSp0my8Uuo28NARtlC4ZXLVRwtBWxRRuM
PpN46hJEEvBN+XIMOpb4NmeOefPm9pnEoGFSeV+NEmEsplXI/UEZxnEHD/VJevDECiWT2n+SZGmz
HyYGkMcE87S9DIgt8lvIZUs9tHWIpeA3VTNI3MV0dn3MM2xTHamQYHIBd3wnxGeukuddtDTJatOx
iixtIdX+KfTvERwm0nOLvZWFSSRnzy+acqXnc+0YbXajhYlONe1E1am2kTwJivCnKBdN4Yjohnlv
I8ivk7xy/I5EpzBdx+iC4JMWXIdxXrYarFeqECU/3PIjgx0RqPuMKOWsltcMrNUQdC+04gPpEnO0
GIwRc255P1UCMDYRuyxMHFtYm2L8m3yM+62x924t8Jx80X64FlMOhvoQV2e0MiE88glegmzc+VnH
ISoHdZu0YazX+BDLWzvSvycXA+Fb+DarwofdRGkaEovKmBqaC4sKL2kzMINOAyxcMd4Ou2qZnE1w
OnVQ4iGNLGwAxTqqSzQPFvI62e1a5kxsx8WDdOf/2oMAHzVz/LEbnXg5gRAmg0k3C/PqeiPN3Yl3
AEF58wSRrtdz9J3s8agObDOqt+1Obrb3ZNMLAbRNLcgBQ1t8sJa0CP645bNqfdLG6GEDZlYNt4ne
XFDD+TODvVxGSwjhj2BvQ3v8H6akKl3ev0iRQC4gO3+m0kKIFyUjCCR5uTPNeRC6jpCDQOjvHk/r
zaXFxUhTm/szuKneL0eZUmLOVxJ3oBnBsPMr3pWSYl56aOPFH2qoCwrNosxdoM9hoFvb8Jvy8eGu
45BxTFjykgvQbXHb53iyi7KyRDoCX6s7AYHpUmAlmGDfZHttTwq1a4eI8n8mdbIaM31fZXRif4A/
TU8k3NKw7fuZX+VfI1r1YjY8PJ2PGPYEgzOmByihGO0tp66WoaXVpD/LYKIo6spblYmuY7/U18W7
CS3DpF9yiDXHRWur3YAX5+zrxXipx1aA9aXn26CRLslru1GkgKre6onVABibRLfzW6feYgPHKn9w
ZtX6s/2VbWWI6k2C7SvbCiOcIp8kiV2IPklGrCoiIXOoyAJ+YErRT3J1zhWe9PZy7dtfWAR4GFMo
qpdwpY1hzSWYnea5C99mbgeF2PdMZHFI0oSV08pG5E1rwB6UPmXO3loC1iVmagbeIcRgz+i5t/j5
iesqmVPqMuldhUMxUoexHRkZHZ8d6hzV9lzjdxnqIH2IULBRIICJE8HnqcrlOhRKFxjhwOc6dq1U
vdvrubxRLhlZJ7sR4Ot3JdfGoGwDJ+eIG2Cnkhd/RCGT+Er/1Uf3Vr+byXSgr71c6v6Vm4Ra4E+x
JAUhatt2x+ZQuZPlKrmWkYOhpMN47jPThJf22w2Wz6uFkxcaquDN/mPKh4IqTxVcYTFMlnFL59ae
z5XZfg1agjbKyn4/7vwJ30Nk4Aiax3d9BIgg+RhQ3rsTRlNb404xSSyC9+6R3ldtKyWk32AKPXot
a2BCOuoZu18GmHoikZSgLWNM453CvMDDecgIKRqlZlOEWi1M8GYQ0Og/uK+MRheymDxliESVL9kM
R48+LgGHGzT/Drs9OHDBkCrzVsrQbYODj1zvfQ4dt6YZj7HnPS3T8ZF0tH/oK6UT7GfB6GFGEQ4w
JztQ8v/HS/8XdogXxsK15eeVCji5K/00FVoNk0RWBEUUe/EWE9iAhOsTTFLkAQ7EDHKO/ccih7xK
xVivLGlh0EFE67X5ths+L3uPoKA1s3l0Xyeosm8qygVDDJZAEmXq0lKXY3h+P6HERMvzG/UFYY3j
s4m3s6HO8JXL8rTurjcSLMsc5xP4e0Ag9WNF7UBT0XkUUDVLzwf4owi/XhQtwEzbrJqHABfIYztK
brHl16H1hus9rdi2J9v8f2Y4YlzGqufU18V6GNQ10UU0g40qv1NqC6RWkRzbzQK6wPBGZaHNGMCx
Y8IHz20p2v9v6KfzNcqqyfMfj67NcpsJIG5BLCPZRY0QBjS6L57V1eHuCaNzp0oC0+8yQ86axr+t
hWMkMqE6BQeoLTwtvPtjUvNLTJd42I7NIvgAvpJZPzQNTczPoimMjVZ5QaAAqMRAswarBU1GDckl
ku4ruVXy3G5iYTdtgqoiL+7zALl9Qi3t5SVP00UU8vE+Cr4Vc3zQykYoVR/1QNO3eUqJyB6J4obl
h4ux+6dTEfskiio2PjdKgYRqenz+NbmR3PoTVpjPoZTLS8WYYzqoy3JFw/1Ua2RYVoFhSSQDIkrS
bVpLsUdNKzjYxshxddX5fLbCqAJOcdle8kgXC9IB7kPuK+O5IbZocGPZOv8TJ6Plbwcmk00HS2Fj
Dp12OyuA7+l8V68LwpmSkWxjD7RrsptT3m59karCLRi5mKYWgFEYU96AB5Ogqvjm8SwIm9ai2tW6
iLfjhTI3ljDT0Gg7Gp64R5btV0FB/qrkNVOMoIK9NwWKig0vcjZIFUVmDcLnDdC2B7EBztRMesCS
yzx+hDooS1Arsrb+8AWxgfsM1zn5cjkieZM+Pi5WDn4F9wvD3LXs7X4a8qJ7srjrRMOkOjCCvxbs
TCBO6PnNzQmKyaC0GP020KWeU+bVtrkei1npjJSMA1YJq0KED72tByjokAVFPT+tF3IPdQGgzjJW
hnusf4jD6Mk7whFLpXQ56cMEJbpiTpONunNOODQ4kmVGzStvVsmikmg2WDaaHV247acSCr6ydamo
i2OOHbaPQsvSsaQ9dSeaxIYfN0ql1xYylKZNGvS/w3+Mk7HPHeyuvrmHvtiJlOhYqDe2k9v2TweZ
fxucI3T/KtHanbNAUeDMkigQE8IwOK3ap46NDrY2CRhDtFU+sLPQYfK9Ragw2B8CmshpqV5rauDt
SOor5LYwHE+Ikmiwm1p4bRuFJTn88fj95dJW6fPY2Nxx/Xp61BHTYypQAfl4hbp5a/CYJ60+6HjY
mDrKO03RBpw+/t/mbqgOlmpVTU+SmLcwHRnxOIGcx/Ej4WXFz93onbm+nzkPuvIX6o2RiYEzzHj0
jFWE4YnWn6NUOtAVQt3xK+XcB4cLZ6ND7QMKG61EXeeH/ChIpIjKm1tipZc5OOsodyXPjVRrcjeS
3pp9mIeNmig+/oUn/ENBFkV1BYZlul8LY/G1c7yJEGIy2z/KRl6NAN8pBr65AETZaYa9p6H/Sp4A
WTFxpmgwszU0yxwpqj6dpvmjO1q6y/CiI/ZqWmckxtwxCPwU0I/Oe3mcYkAwXtjbVbs++ghYBIFV
iYO0fGrqGOfFRQYKqhere6PHayWRzoPnjbrSswLJATgf6CHkll6Hbrmn7RAi8iyW5QWDv77JJfOK
dwdF1Xx6XbGpvuMznuWqedEhs1NQQd+QUBFUDYsWL8oEyWDkVoEUqPvKVfcTUfLBUWtqggcoy8QK
tAgdX+4Jl/V4VPvdPXhFSZf93HcYUSqw+bCbf24mK+sEznZwmQXRLvQKOFM2OmHdle3zSx2rDreH
RT06scclqV64GqU7B7OwD+9cmTuty7ZBnVraepq84hMyh7EmOLvxeAeFKOfzAopSGV6RamWb4lYF
YknWpfhhWqQmlMJeOZQbgigbBnD1vr7qRmUJMfggxdUdFEaAJXIkCbYDm9b0DG4+Ro0gTQYyQQ9N
Hmhrpd7ZFyN3zqG8kEkj7RvQjwNl2KMUZSiBGzzIB+N8ImdvynfbtjFW0HXA1tnPe10eYtXmKqmD
9/+N++tSAgHZ9qYv7TEtVJpgCy5IJqjdhBrtkSTPe0Q0NhrQcYkRS5tur0tXfYp68V87nUJyRtcN
UyX8XI6akqZnjOv7+DU3d15G5fAAGQPfPDuvMfgJgQw0WYIKC7Otfj5au58YJ8tUvTBDEJH4QuF+
6TFgTch+Qj7ma8bIuEJdJ+CaosiHVtygr9xQOogLbPOKbbLG/vL9NhOyCvdz9i13pzGeVBcIkcKe
WKAK1Rihf5j5PgPmWMhChX89NEoNnpBbMR2+wIoIlD0msal4yB18d+Xox0lyq9j7llZgx3/8elEm
VNTW7rwMonkkejHd+7LGjulTMI9Ihn01eaTL7GzoW7XEcQ+vnnvPQk8UsfuW3ifPVAg8AXPIwkkv
8+444itEkJx5oSfE2/b1EFE3630WRWxKVNJUT/hO90SINxzvkiVu0V6L2cSoVb7zZmnBTT6lzqjx
yqprsYkYztMUmtxAhy1Gdzt36iGFonqZ3YQf8wRLcWqIm065TGXhUn4H/ePLOKFsCIqrRJBkR5c+
PkT7ZNYQ7CJj+osaqUGGJXTrq0Cp48zPh9e6j5DbU+79sE/QyER9NSD5OPOC+N21FldaMRK9wyvG
2JRKMyoW0ffnV5a7mw8btQhj63BCNQp/601zKJqh8vmup3JOFb14IC18Mlj0DlHMqq6Moztc/BPq
bkHNXdv/4i9wWzuehjUDE+wR5Zdz++8RkKcfK7XkO9UeGD4e3SW3jZhK33yxzKv/Bz4ikRptpxW/
T9JWoxDHqxtM0WzvH2FUoH//8hcVvap9am6t1c7WRHwOWVgBmR5nDiVDY2oWMbF9YsUR9JxcYDuy
tC3n4vd39lvEJcf4Vw3SbB1hJTW4lMc+toj4EuqIioT8H1CN03F8uDDOHO6bbSPUBPVg0SEKha80
TLRtPo2EejtgCJ1T15W5g/nSTHxCSFZpgWaGYLlP8izkTzuW44QImmKeRSXb3DftmUzYfbDI6X4l
m5gyFqfjc3XzzaFuielRm7kWPnTw6TQTrlUGZx9b39Ed/amWCjUoNVCKawjV1RDnKc0nniSB2doD
wS6ZFOtDMYlCqc+uC8uu4bKgReYbKoEltqLQhkpbWrvclv/4tKsjg52dK1vxMrYn0NnNdu2mbeDN
ld4ajrG7a/90G4sAvo01pceYbHkbixag0O7AKoqn/AdXFw/85KHoZ/uRLRG1kaLYftODURPulDd6
vBGitPgkTzajMg0Q5sDY8JxUxvYQXkK02G5b1tC1Cj/VNl93azb3IkRxLqEN74R9yunmjGFi5EQZ
LxR8cQUcUPW62AqbE3dJ/AD+PRSpzZkYyh0FkJcSl9nwlPijPxb9GkjxDouQDRTTj8AJjpEKyKPa
DJXbJI45OeZwnJloEHjJoJYm5NQGRJTxNIAM10NP/llMFVW+E9q/++xGTXj7poMFRHdAwNpvoFYb
uCJuUEZ+B2AQf63m36cJu4oImPbSPsqseAv5evrPEsCc/pg97WMNwDV5cQ9Teklq8d6/sL93BiTI
eHYyzvZEOzVxP/pili8L6f6vM5yW7qik2KAjzZdzCdpgbaOqLkJTtNwcV4wLZnOgqwLiYBv4v4my
vQWKv7brlux+RH8/BEeHgFC/kYbJeH0b2uUlXtY5yXy532acuIXbQH3CoLr8HYZqn4zSC2Ykr4EV
LG8T/nX052ZOUPblsESw2Hav1KjQWGY7Kxjfy9O2mscZABNGM4POxG/TQFUHo7N06BcfVD4t93gZ
1qZONcKPh+8WnyaTj4xNABQOVNty7UNXfxbTVsIWkCTMKNnvnsIzHGtTTg98gFaM05jjm0c5e3rL
MIADNWrOXzsutQ1hJE8sY8eg5qkv20nvi1lP+IdoSYcidYiI63VimrzrMWeOk7VnU3e7BPUsnMFR
D0SOLUYsUb9Xy3m9+AbJxSAcOwbMTCE+e/+HauuGV5eZ0kxBEIaTB2+CaOsPGZJs0DTOlueXDnha
rQn5uOnr2LpCUcmxgeOrX3oTGjxRp/1OUvwivETtJSmg8jdtohl15cuGql+ePRw76d8D+9LQg4of
NiZcGizgvcBE4K2ZtGMw/0h5o+gOf9gH+bsEwSBPRCcMfIYFDhxRMw509eu/P2mYUhRbmlqMTjjL
QjXgVkSdAupP9zvNGWh88nlXr2fxVYUO/oFhNVLfA/xJ6+sqAyLarS1FzmmGXkUMmHFil5zlfBjl
treviDy7n8rsJUSNjKK7AP52TG09Y5XUpv/2JJ9Of1trNvtzmc2TMIsmgEblR0/wXw4sNfCjqc5l
WbR7vf/WW/bXnjmEO4Y6aRrXlveDmSDChan7TAC62C6no/OYv4Ivx77ZO3s57wkIOV0aEuiH71KD
1N5+fUoRbG1RDLxr2vK2khnCO7IOZ0LGmTHVa+rXNKDjobchfarDVdYticI/CQcomvsFMZtN7uJC
8yTygu06laXcUlV+wIzpldZ1f7Jmehpa1w24FS40GhbnqFvW7pRI1IhoC33Qr1N6QYcqt6146QWq
ffBo7KJIp33tZWj1Cln/2dFmpclGdAyJ1iwRrY4wKtvBC4gL5tjAoAmOCXUZkD0lLjTAdNBFPwjo
ryskpbNDrDy/Aq11eaqwCxtKGlubnmx2LFpnCEMv9t29EU7Rk3cwutpBRjtRJyxx6X3fvDjoB69R
64bAbaJpi+e6qKUt9X45RJyx9sFg4Vuuj9wJIKQJWwZ2d7hHw6Qb5/HPf7uKNQfGlkCvUaMjMHSc
ZOLIAEGjMKaCUkK0QAPWIa62aFgArBqsMEnfI1v0/6i3evinUoML4gAmTYh0fc2tyMeucaBRM1B/
GZu2l7/E97jKp1c9owFdPqZxnGQOXlnH5j6I5naqm+rHm0j9ZrXlvBbUedDwHqzRTjUG3KSKU2Y3
LauIVJq+N1SpgqDmm8OKr5I9elKO5uEVOyvLz9KluDHLC/i6mBB/rl0ioyuTgTq35tC9Ej/1q+XG
SqQ1w5LsQhNWzTxzUg0dMMUndmPWcx84aZvX+mUsHgoYutnY6fvWWEBxbJVcsrqwkd1ucnc+uIhQ
/zQQGZCXko3XFT4XeeW4LAZI10Vy475cZeb8RoVSTU82/i4NQ9374of0qQKuIOgtsdUuiu0DnhpY
/cRVvBTVQhAagejSvWfWW+PY8qepRAHblEp19o76oicXOWzPqujbO3gxcGmqp3iF/i7AOaUgeJJu
NN+HT9T0WroNZ4MHOuUEHfVOLH0M19zNrbm/LCP/ThJ2pRNflsH9kRTHIHCBkFGrsa6bCkzo1yI4
U7t/Orn8XcoOpjBI0yuSVDH5EBfHUXVsfpX3tUwEb/j/LoK7qjy3dkRVamtiXhptopVKEReDIaHl
LhS2fYPQENTXGRTrINSK1sFajjXmYYrNtQa0x7eldkn/k6JROcSPkAFVoSGP/gizw5YNSae6LVQn
6b8IvLkB+mbQLI69MdwJOyRuPVy1R3GsUJ2r4cLE+rK6UpzOGRi6bkRWTziyC3lFt6O232D8rcHD
Io7BStM1B2LnwFquy5c5BK91aT6CXvP/0jR/uXGirAAuOg0gG3gpIQVNPVx/5LunYAL5CM/VSXjy
tYoPebVmW8/qWDW355nV9JHMD+igo1vO84ETppFF3nVopmYpsv19BXOs52nXHnyasJov3llxx2MO
nwvMjPLy3bKiyREEgerANpvAeyVGZYSGz/eSiDF5nI5spRSlXPryQ4h4TQEkpyW0QKWehWWYfReS
DUQx+AzLMztdCKcha2y9gojY4JJNbNbOEAbsSRCulInAXYb4f06Arz5a4+c/huPxIdbfDuAkk55m
wLfCGVn9xCNV+yesx0/xTAIxKNreIkV6KrC5+mI2wso677y3ROD9Hdxpe7kqauxaVNg7eyPPluS+
edZEqmsdQnpF8UtxIW70lNAmvULkBdBzdRplYNOBZ8Xc10QHTdlG5oZBUne7VPCYZHsLxyZFHsIw
dmk7xzRGrS0fTcMF9p1jT2Ko+VeyMiAd0h6J81Ugqs1H1rO6D7O+xYe7se6nZeScx1fAHJYs6rTD
JlzSJYtzHr03CorC8FtHIksR6em//NERafPLMIOiF7HiZXaVPXosXFSvX7AUAoWkZaWukH6UIOxu
Fmp4rrbTLpG/I96QHdrqifLhjHU0waIo5krreXPU/L2ok5jpZug1xD076NOf8wJbdG1ueFdHFt6N
W25zlYf6T0kZl3HOIj3Vx4mRjO4orYHH5von4Z4BCsYZAfNtCB/FBkxRTk18Z8r5Bx+nxmp+D6Nv
Te8fbOB4KTST6JmZVmBYr/ptLqRcDJ+xu+O+R6t5sA9kSrAs1p/7E2Jhw4OFuuZUBr/ldqBn1g7P
UijXY6+OW425AyWm0YR+DbmlIHDGX0VBvuR9v592SYy3EeDH3h5WtMj+R4MmTgOW3+Y2x30CtYjo
6AMVUthEqFBSOCM1Vz3wzVhIDyHBxzI2GvbVw4v4sacH+UjgnvRy3UciW3B27thzNrQuNPZ+ifhK
Ey2hdQydFTmO1j3tvmVItEUKSevqy6IRYCCjqoNlvInIBX3gF3dPf7cWYzJTAG97TGo9/mKnwLBk
V559P6VxXzA/3ZMW2/VuxASOJgm/IXExhXAMmUSmcsNaZdNDaqJpwGdn/RqfCFr3wuEqKhOD+TDq
fIumqhORI882dph0MJON2Dsw1VnOFszJ8mdcKU/0kI0blCVBd1RhXFCYsFPCMn0WWYTTiuKiXnzi
qaWT7Wvc/CX1B/ZEOHmlog/hMz+i9MYvRnhZRZvXDU7fyuPXoctjKVblUqHC3zFaZgHuM1nIFeQR
PP3eKf0SbOFc/3umeqm1DP1MADuwMK+C4GYGiDEv8Svyq/jUKyOLQZNQraADxZ4F5Bor7ymcBW7J
tV4QqIhT8/eqFj0q+WzqcX3fofaxMzVHP4NW6XHyockg+RjpM/yU0lv9AXyHRX/QNAsJM5pLB6uR
HF5WMV/uT7roDOH6b3+X9kiMbXRyvlNW5pWy4Nlr3C5qt/bMaXL3SM3p8/XvIe4O0wdOEgUxkvNQ
my9k62BUOxUC4jxm/hxNAbaABiVA/qP8b5BzYgz2/AU+DWyGzjRGAHLs4cQVjM17WqhJb8xqEtFA
iYU5fDWBhCxTjhm2cqjs/HY3rSZSzGp1x10nkAC1n08B/mBBKnR5HV0qP1pHpgqz/6BvlmOu0CqP
iX8SNW9zmr+vJQUtwaX//EKXS5VubdYu6pU+l256TEuOIuV+ac+d0ovlhrO2o6RwInPfjSLpsGYw
jcjnlLWvkgRceDKw6jvk/0zES/u27M2IzVcrk5tTAgdVeIvB89KhitqXsVb83m7DVvIkN5DDFfSp
hjoIdq6/CJSIiIVZ5BTOASXrbXJP2XUzUHdsl+mAnJKc0NRUWhauG4E4oY4vqcJilx5s8p7sDHqd
8uKXnJ4FeAEgCam6l4URfHmWBqCriXusr9KODJg4DrjCwCt2vmnFBW5PzarbAH44zCuwtS8hTz6F
tEVs6AzXkh4teVO0vb7+Yq48Zrho9ktDJI5dPCVUCw/76epC15a83f4y51fpJPE4TgmrzFn/v3s/
QUMQ64fvfN7kb9rj+KRO9V861AD1KwlXEPzQWJPiK8hvRAM7dZIn57yPSNw+e4/HWWaHhd+Zd1d0
vYxH3dYyA0Ri7UQElvw0uMQCvvtFqPAXTTRStO8vwM/iRJVtuKs8xAVYZn2F0a7UKWaz0mNfAQZS
Q+loX2g9Le9uggGd5a2Rz/3ecZIRVBd471UB5XABcBViM4JdkzmRhBHixU+g0w/AsxNfW996qIa3
eQygo+5wicEZ96oSXibW2z9FF+ct6cwMtQXoZvbvoJsAVOFzNwOjQuPv/yDRUEtIsnXJlYHDwxjp
JrK69pvqbzqyHRlgksh6H9C5nRpxl88DlOcdQybRL4PatoCxmsjALDLqgrXpN7PgHZtHTppVnux9
0quyrJpItiTRkza+BuXo7RfZg6ywSTSSAl1kIG86oPWkPLlukC2yF0LXtdUZK4cQzpBq4wtxJD3Q
3qmHBJNURKh9VzlRudvDQeHW3mBcEnYrTxB0eRW9UcuT6DvuKJxD9wRGm4CPB+QQ77Fg+Z+2ZHNw
v4LX3NKtzbKlTcb3fUxKmxfG0pS74k2obkHk8yACSr98K0BqcQ3KJuCRUGRNlseU2EMq09qtClUP
CYGPpjB3kpPmibdgV/MAv/A1dHc/gUJAxTak8Nl6YWZrI5soByUUr7X9fFtImBB0pU7K4WegZaK2
guke5Braip4uG9QvAjCjzD2JDL9aljwONYr9vwLtGmWuzwZQkrBWz86f0qEPd5EX2eZtSyUQqMC6
IfoRxy+Y31DnCXUepKwAw0gT3BlkTi0tropnJ1Dwix62oI67E2eLRuYbWkbsG5SvclSbN3TYqnfw
wdcw+jTR2RR4wSjBH2YvyiwH2tI6/RduplhlyNggrJI7wagU4r4lV6Tbb0JMzanr8zh6jVhAFhoT
R4r9O+YWNKthORBTS2y1T6gUtcCSmkYMFtLEHKRl6ptu3BW8YdQotAHOHJhdR4OR6BsLdZ3i+gVa
AjmlzKQe6vuOmCaByMQnJcp5v0yQ/DvDNN1X+Icaqrx7yQgR6/K6FKxBh8RGEe7bOq22ehDN+vhy
rdNk3vaaeWWqu0AMlS40kFQbdxEgdc4Q/CPNZyNE5VfqsupqJvB4vJLviqeh/y/HXbMRRJEfpQDs
y2jWivHYenqPqLr6KitXs+l1+tvY/P29EKFESWfVZiLXbwyr0qaeDGFlSRq+f/cLbpH5xjhHJPcd
kMefxaEMfz66/V9ZOjsjMMUIw0EXCNy1+kqGrn2epJ+0qst5bRpOh3PWhpl52odYNIug3pULFKY9
kGBej2nH6/PkEZuADGWqJLh20gGKs9MwVN8JZOZcaB6HBCAcaI2CU4NJex0R5HmSKCcUAcV1wtFA
uzsyzl6+lQztI1bVDXxg5/hCGrtC5aX7buNqNGsPTnJD05FxxfWPnDZIafoC7JkGIYfDVqA3Rzni
ct8jry05tDczfGG+uO13wIkJ6OZ87E0tflYplMignOY9LnFMs0I1PGCT8FJvot/Y0j1+ktJMRezt
Axs54X9Zurr6WaPNxBibaZpkYkJZ5ahogMCRqGWMet96vSkuDpSL0xXaLNYuSLgcgqeGIhElGCbO
ESjEEWZRDpGOLO/tWkPdAQKT1ixEtDuC34+0/0nHnJBS3rgOg49gjgkGIyDdOlIglD6ZFL0iVs6M
Vn9s2/kzMaj1ykTGM3G1otTVq2EtxjetTn4kSZEVUPL/1qadTHttt9DjBSsDEG7AkYOJWx6Cvrfy
8QJBycdk5+umUmLs7Wwflm+LmZ5RXVmtKudtc5bf03jk7aHlEM4Iy02eO2m1pM/vhluIX34khzd1
4UGn5xQffj8CegDn9SU/XjODM/F+ZdKQvqz77ugEV+wUuyvyvjIx9ChSjl53LIp3+gDUX/HRiYqC
ep22HZMTAIqVVlAKkBQz+6mW19b3qAhr3NZ1TjxIh4wV1uyTIVKhjd4pK4mGQWP9y9IIDai26eun
Nim65/FJZ2L0A191zsxPAbeECklww3+L4VpX/METK/TSuATvXyi228+LD9tCXDsPAT1RXBJ8y16/
ZoGwqL2aTERa9Y3U1yeAwntbqxv6O539XaG5dKXiTBG7u3jQ/IA0bhoH745HvNSUFKvinCb0G87e
6fjjqTMRn2MEj442bTi8B/jcloLhkBzcQawxCA5a7i/3S0X5bu8sAr9CFSds3wGTdtjENI/Fq3bK
tEGfpJiLliNO5mS4RT3YiUCBkrj380v06skYq7uPavbyrmVrmvhkMWtmGyuQjzhclxUPvTaOMKaa
qI1g/cw7c+Gl+J+wNt7v9kXV5dJFgkf5GRhh42kypUraIS+3S7xA+qqQJikYJQw7lFBWl647/kdM
3KdRkrabrhbhe9VoIgysLY2lm5QT5CvZmqyh+r2ybkEG/R4cgY1AzI9R4xgXT+rQLOdmiFTRgpWh
YnMuNdemyqNrqHrz2drIe2emc8gcmkIkjI5liN/xOMhusJHjF6OvMCQ34W8J0fuR+TYLRiQGhPF+
mnX8n9/v2tAq48aL0bc3lnSycpYwXAYxrO3KB2qDgK0hXsY5WXWYviRpYC3Z1nkJc6itn1dERnR2
cE/8+f3stoLWc7MeCtWUXYLB+NoUIVLmN9AP91XpvvgfcuaB62gjna7/eERRlK+4BQzTd9BZe44u
xohsm4FQXWYq5VBn/n5Eq/8MAcfok5bVOyHXal28jdxmHNMLRZUiiuLUJyqC0q/mOeoHAYSYakye
z3BXbNIKno7dJ4W8171P9spErJsnXS1ZMX3f095CtECSn/E3bE7/HONsmmi6zs5NPzU1VqR9HPct
7nm/+0euhiT8lzcoqUxwY2VXC+I+fbQjDcRiWRsjl84oDt9u0fC93Wb9BgqLpEKpQq8C44CRs6CK
OJ6SZXxjCq4U/dwvTr7TN82IAl4JBMUvd6W0pkC6BWviNK5IMIP7WH87gO5LUKSpJ4Q91ByMZtCE
uyW7OOVYXqOUdATXQYqco9jxyZFVLzgd00PywMT0S8lE5WSLL1B9f0mjRcPMdIOlAdalS+aMGcRB
88MsM3xCLPK0LmGherdmjJqHiyOEIZhY9MhSBV5gtE38mG561ABEACP/UxPWUpLYcwqZUAob5t6s
Me4tNM9khdJQIPVkwsiZph8W3ET0mrNf++ahdxnAWlvbJVCnJ2vwtvXSFMIfpIqih6OONTAEqik1
SlS3lIQbWxylPiNDjaFBho3RJln2JIWs/9i/q1zoMzQE7BSQpa/vDU8A/UxzrlcY0tapB/vR7h9k
479k5KTURddKBHM5Op95L0RiJ9QqQKEdmPo33w9GL6KJkcfsnevZmkl2w7asP6fcgma/YJEDGksq
SPYyjQ30TVPxC7qDmbW875hIs76E+zWZFPG9kgLDOoG0URCBbbSMAZWEUonkiOm42f9E2ANlEGAZ
WDw4pcbqv50m2/AExtK5pO8GPnTdvKPcvN/T4ocAuAm9gUQGWNnGirRx7GFf2Cb9r/xkYtZnuK3T
12jrkuklPVkm5qjNNMBsQ4qup6NbxiFVk5pL2S00tsAdInRAAteEFhGaOPc68+NURuwSYNu1D+6t
ZgOq2f1FSGnAjGTWrXgRYovdfbxZNC1gJAL7guVqMvl4Q5gU7Es4VThBdH1XufmkHWsiBKLQbcCA
rUkgaFvQAF5TVUf/0fRzf07nl6Cubr/j5zQQp8yazGYrbZYoJgelkxeKFExnK9rU0CC+uEKQrNZQ
oF/WHP9XhM1jIlsZPdHAEvGSXF0howNAs/4skvDedFC9n/Vtr5OugvOiBXbXPi/X7SJIZ84Q/RbG
XmsjJic9TJHT8lcVMF4Mr0vbk7JAv79J8zJw/LX7UFnn/lq+yPFIAv3gM0vDk0QmouKgwxQwHjt4
bPe5XXw+AeJ2aGFWTpA8BeF4R1zY+W/SNn208XmWQpec6cf6bSDBVZ5a9tYjynZ06e1rZwgR+tU/
Z6di096iQyFtmjyFjsRre8EDO5Af5K/l5cQ1X7MRfob4cuVlNb965m4KCqfh5CD2kVxNWoFGI4bS
5rp39rb5fephvLUcnZaQr/hVy+QghDph4POBaG+YC1igawuQePbelPuebDwCvJHPMKXwqOqEuqPj
f2DJwTsN1xBBA8cXaN78BCTKx4kntxjGJbfnOoE9gdd5mnl09gsPkD7E5PQRrhTf7TFF5uMDfh+U
YvgIKR5sEGhTDAz3J8WX8CATioh9mPen5s9/jm9N6kKMe5K1G0qzEyrgAzh988QZ3TlI+2ZbOxM2
N5R+iIMzLV3HtUSvQYm+Y4p2KeyW6qZzMpMenLWRNSodSEYavePuPp6UfmzBbVsJZfyB8lmIW2qk
X9OYyiptJz9ZtN5oLI9Um128N7wG/qcWfRFtdndKcNQz8brtEZOE0a2gHARlNtNFHOdKpDmMlN5M
97ClLY6VsqRfpB9UZPMhlMsfYHESDLLQz8VUHI403LcdjJr9ofUI/VBzgEpCpJ4P7mjMu4cTA5uQ
9QOMcysMD6mEhlAJ/51OyFtADs0v7ABCkJLQXI9H3390sOJZFmnb1dk4cmxgS1V+7A/AfMORczyb
6cEuhTFwWTesdBRgncvpNIUMXEWiTSOtGNrGt6WjrZE+O3iqR9jpyz2MqxcyblxZMjqdbw3QfGyd
M2d3DFwems68Z+cGhR131xfz3PQKcYe13XeAFWtB98sm1DLaDvva6PQqyZ4Gw1d3ACE4yWaPooC9
9eu0S0zU4XhYa3z8KvlUo5wI2YkD1sBb6PYj2vEzVa+OX2a5AnMZrUamCj6Oy3+5aQevOarcgCNS
GVmHoPJag1uhtzq4z7rgF1YsUGEUNDbGXii1MUHkdnqJWM7bhdiQu2YOyxU+QAJOkK65JsiZOUvp
kzIDeb1UNAatUdsIE4FwsbEgbWZEI4VRsPdTXwTEF678Zfu368tVJBv8Anxmf2zcfiuPmYh+25jQ
5YThlc9z8ZtgleFjaddZtGe+VYMoaGKxoO/Kyqx8CDvxdXzYXuuVmYYgy90KZRwrWVwxL20+ABgM
sx/8VHTVejvytpJzz0rUNLdXChzlDmj/Pstb0aK1ncfqqhdINKZt1A2z+fnxpSccrQ7DKTOc1vVP
fqUWl3be4OSS36qOEN7KIt91PRe7I1L+7HkjYVe4ssAnoDBbVy8qBHwdvNJHmXw8GgS662KjltsG
2jVyIbjTafrPX2MkyNFunyjhg26STG+2z4cRCWjfs9FeXHUlY99vpFGb3/oXuAHe6DWGaj829jE7
ox+0D2jhFg/FAjQow8+Kjw65GyMzkQorv5t9GOGrt/5YRIXlbQvAe20c40RLr+d1SMN8iQBr+Fm2
Bd/Kd17qvbaRGIFjXeNqeHUMtVzCDVYhJupkEpQ+Hdi60dDkP1PzfGzWou1+GzAkrQCdrCWj2NeO
1JgeIgaXQ/wyfQAfBEcsem9I2xl8jduYqTgtXGzBrumSZJnUsJvm+bnDhDXtT8KTnCwyYjIQijBv
zVGNwukNzoz3pK5+OeSRAI2PMjzBHEcKfbnnBbFrASc2hoRzBsxtPvJO/WbNC2fdTDchX9g8cLhP
jF20BtwbglplSplVpTDQb0DNpDKHyokzK2a71NeRiLnwdCiHOju/k+i0Wipx70c54V28Dp01KENf
il9tSsUqmw1EbsgCSftqcfno8a1JBoDWcPAvMD13f3chTH+IlVPhPn+jLnEzbM1wY/a2z4CZKTMU
xXbIU6K9fJ2FA8l9DBpJJJO3RLBP+kp+UMPmD5dUbHWA3zRIlamZSmgstyGPLGlNzI+vPLVzqw1o
0/1ZBIfTvEVPLeug8PYez28BWFGUf1MHITo1bFuCrJim/miuD16Coyn4haEoCIQZNuKvNXqMYgwi
qXLijKUbf9NCITkoGFPAz5GD5e2aJCDgg5fmAoaHhqSlDz/tytJaf8Zhuq04XkLBrGMqFqFdpcDr
L4pLjpQOmrh1B1mS2s1pJQlbU7Va4IGQdHKLi2O1eUQNcfraSq+91yxDqzeztwJe2T2b6C/CJ1Oc
adS7KQ7/cnPV8fgGVp2bmRaK3ZGnGwPXIuFIdyTopS5uB3YD2RSRc8xMHFpslks95/l84yDrf+IS
hvDKQtyVS5jxxPSz88c5lPjfmXLDcWquhXYBPBlHWaVYHzFxiMNEghfsoaihN8uL0xngaBUvc1/T
IK3i+H7YYfMx4mvuGH1D+nVrkvNDUNfLZ+r1p0ls4EBWPRB0L4IAWKgCIQX8MZw2sFylQ/bhAM+a
i+OD9YDwTdQGV05WBKTUohkZMrYOlJa7Kws/1vQViOWxGJCCWNT9r+Uqeah7mUo6LcpSH8MyQpL3
gKzYmDl+lPxrh9ny0O3d/VqkiTFUvf1glixazW1vHHCQIBsqmL8Gmm6IDGbrLJh+bdPxurfgK4pl
00ekcdpRo6N91vPKuBWSuwj2PBzYczSUt5SrO3R1fVtU1SBYNAFlic6Sb3pWLkfwq9JfFwf6vKRO
XtQaBwkrsRRIVXHtzIODX+2PvavHxP84kDWbyn8BAsogIONmoVLG+bUoYdHgEcvyCU1190HyHJoF
A8B7y8m75tFwG5jIoQJxIT4IKqEGIYGCrQjycQZjPobSyrl34dQuPzmcC3sDs68zmTUHFTgsD2p/
OmDN6E12XBNWLgWCFIPilQzSAnV9+bHPI20lsq0ARl34zf+SfmUvfx4bco+vgDjd9bh1bDphf9T7
zjWPUNqfmBKY/fR4yu1ISYFlfS4ypJs5SVNDCQmtAkeWUVjrWb/suIs64Nl2btDMJh52Wni87pId
K2hSNGCMa/dyEytpKjkdp4ycY+4J0F6koDKDloaFj9qK3j2Pql9OWflZ/vJ3Yuqz4u8wySKvaCDS
Jt2dy6mopCAuKNpuRNELW6r1boJqTibQnFIQ4RosUQR62SOGZB70DcV/4b6CrPhxX4wf6CdDSkWi
qvAc4m8c/gdp1aKVEiElU/c7ai4v9xE0yrw8qhe/9BfumIEson/EigIFMaNAqbr8gQOqj7+gddJs
9mc+qy17h4qo/MvVjoRNf43R1CUbIA9XqSjGiPHy+/Eb2bNQof8rnwCS+vt6tx5cKwIhmHJsa6ah
dKBSDYmH6hPaYMuVlqOI52CeQJ98E9kjDpGzwOisqJOF+FeCroO4/ZO7mAUWS+JzoJfcDAD1rfwD
5utKMVna4YZKEe0/U5iwWTRWtrTO3JlpKR8VDDcwYee3JZqrm6p33J7qtNxmVASGZl1rBUsPVFUt
cBau7OK55jN1Z2S6AdpgOMtKEFD4Z8B5Kp2bc96rpuQRaim04q87AGZ0h0kiHtnGRkualxTBczqT
O9njxOT+W0HyLNm+0yg/jMunGhDz+pw/3IPL1VgFQfFRqQ7eC7Ij2WDBT5fYHBAlE7MCfxEo56uV
eyng+nqGHzvmbAKzt1FL7fvlDeCKVC3rmo/8ZQAhs6jPqvssO+/7Jct7w6NQ+oK8dsHYmBj5aMLR
NZtqtEMTwo5/KZV1ubz0lCErWt8A3qPbOYrbwzadvKxDVb4kmJf5qSM1cdfbhLc5MsDqs1/lZ/m4
27bs70ZuRSrkfdJLjOeI3ytplm4uNXZYbcx+QuSehN5VjCd4/2LEYUu26YBwG3ShGA/o1mQhTd40
zGIestKLtYZ8uQlmhikxJd8oq88CIlpQK80SEvC5SMKwvMTZVdJCwOSfe4PxJhjCB7Kka01amn7D
3zEYV0S9pPO9vhgqHoanRDK8B6Ghv/9TN0yI3pl+PhMkwjbyK82P1O0+ICzt7lZrqeIFcW2SWW5N
PgsHCADzaBXb6/AziWaMQ1X7FnokABLg29GWB0JM6pG82udrkrRQk28f9qc5Fh8ZphNR9F8Txcqk
jBhJUDnFf7IUw4ijbG2gRC6VwdmjVBuU/WwcbSekII2tZmjdlkRFWbU73stQ/TUMUlxSNH+fLqAO
5SdvdPvpkkxQlg56Hv+R0zAVs34QVKVDvzOez7wnRanH6VR8PBdfBoSYR5bT/2lohfFWixlMBfAN
K3Tr5j5bo8/GQc6H9wphfR4tssEXp+vwbK1B3UTd4bEd6kU8HdO+nM1ZQxBXh93x6TZH8hXG1Pd6
HPDVp+Lb1gytfWNb2T8rGJG7co11JPgO2EBlLGl6GLbOfIG1rxYhqLLMqAXUouPNy0saJGK8nojB
sJqAPHs4q+9ME3Yggk8DschBxO430csZDOAb/l9GVflEuUBU7otKpl5rRQ5+1bWgj0FNUi0kRYKG
Y46RWXtSkGH2V8pM2Hq+1jiyjuLCsqsjcn6WN72YDu+MkFYT15j85RCBVGESGEo+IH4f2jtkHaTS
YQZR9kmsxi+TG4uNA8Y+4GpqWXfUJX+RZnkO2nr1zVbggxbfPbHH7rLRydlCAu16j4BlJDVMZWic
q/fAKNgSx9AeSwqJQTlHqcVPoLz7+HEB4iX4wJeTtKAIuNBKsFZoUgPw2/7cRPD9CC6FRAc67b6z
xJBAjbjMXzMT9I72iHSI5ZK1/xU+OHoomNfhtI/uaDH4n+itcITMh5cmREA3ecCn/lWgkh4UMD7N
2DmaOqOc2neaYraw0kCZkuU014eJdFmeKW43D17xExW94rUJD4wA3BZ0dNtMfocU5u1VgYt++vRO
LUqMplc2WS8rGfMgFAAwjzZaMCMVIeYoEWWMYwx0lOK6CYRludS+TuKy/gv2VgEBB7J0FDFYaTmO
FFN4aSZ3PFPWXvYETRHkrFTnsU2CilqMjzxuXW4U8fcZGf9OMW0BGzmVUfewcJZzycmkkGaIzTgg
Q9LgFYE2t3fjhZoIxL2wW0gwqfMxXevU3TfHRFCwgXlkq2cqNPBWErU/W8yxGBkknOfKNDHpuIgU
r3Yl+KeOYX0nysjLUsKpW/DxymO9XOpPAIBne+ooCixrH/kuYUtLJ3obEkvlPq68Uyvd8fogI7GM
9gzUi+Fr+mDJoWrovT2OjfA0j0uOpKx8isXeQF7HxFS3ktfg535/i8FcW/3wXN5FxJcfICWvBSMI
9LIjkUHvjlfjTcXttQxXJ9jwlm2xMg5ho9MbbI2y806HnDOqzEB8NHR8kcm/B1ixujVkJ7kVfQfP
/6jz6eBYoVsvtVxOkRZlgN2PJG+ylkaYKI6aepanA1/TsxdXgJVGzVkBVp9GBkCWZxUf+YdQ1NAJ
oZzZB7GIrc/K7dL3y9HtiQw8tzZfvP8Q67l+rw9K8b+6B/hNPRrCdRYnOVxsxt1oLIIdVlpQ4gH6
J/FNU+6qpmTVRtvPZXRhqHpitsieyFcDIcvzelaGDDwOCkzq+Kv6QkunOoa4DPzM6XRE5zkY9YvM
QZld5ildGtt1HGbu2IpLp7hYtCmFkR4G9LISMto2HLeTGE0sLCaeQU9+beRwSkuAQ/7EjtnKq095
n6JiQ+ft1d0GTahcQEzeVwcEXKlnVWKyueN/5MRrzcpt3GTh16hwTCI9JWLhEWdURbvpEpQL34LC
LpTJfiHu7V+5CEEVUxQYFkkHqaTVM2USVFYRtmkcIWRFH7asenNy6QOqPASfektWVRzyDNvI2inT
mRrzIS3XljHTBFax5iYtAAF8za7AGaffV43I14rOwRQ2+TJyGk2biKCVzNuhpUJDuqYmsEJNPWr2
lmUzmj2ZytgLBClFA6vngaiHWss5y45QSqQXeqYdPEkR5Af9QZBHoUv0ws5mTpdqMdTIbOPVBmVA
aoeEWp0Y736+R9RtWs1dD16wwyFi76Iml8HycBalAlFbHfVq5hT6w6KL1cNvqtFkumZU/WUyuMGk
aNRndqWmMi6tWqTG206dJfhWRETr3InVy0EDy7RSfMyQiqT5SaFO7LA9/cgbVfqIDbpELs3Km8I1
zc7zN1XTPFUxT0hr0FJaoIyrj6aE006KbYjDv5bEwuu9h9NFuLekjpxgnoTRzqgsk+ZSwoizzTRV
ctKcnb8Iza6TE2+LBoGEJH9W84gyMdqHbWEpy2Y+Igbqj9MJUSDX4SDC8zeEE7KErUFrqMQ3M84A
kSmKU0aNC8IAx4+grNTJXRJp6kyNJdShMoqoyfRdjIWI00iSEjnTYxC6VrJHH7o+t3Cpf/29v8/x
y/CQPZU75CbQ4sxuJFsfeU2xsD6w2mN4gZ8e8FWR2klAiJSbFAxYxINcdfAdSx6HuhCLZQ1a94sy
0e3pe+EEIooyBa0kwuFHn5KB8kBaNwlv7HZl85IFGOzfRiJIv310GNs67DqAOLf8bNnUdMPid/20
+062ZZXAghn1J6jHXSY5zP+scvZOUD7b3pdhUfzCWdwSZ8Qz+3rj+bxG7dHj2h4hkU60YUU9SiKA
r/hNP83w47+Wjmu3Q1Z23GZR7lGWBrSklOnms9w0w1CpmmZWIH4/p2+1lavEuvo8WpgLpuCrwacJ
BF+CCk6Bnw2k9n1AnX1IE7KtLBtmkCfm87WyIDXocMjPVpW2kLCr9XSqkRxfjJjnQNUmeUWYQm3A
RzWMEsuocnzFUuAuGCCZys6DCKMqOmnP1pVbnH+9ZdvB9bUymqXITgy3M8zOYtL+1oYvf/zvjPUR
jTGYTPz7Wrz7SsmtQog7gDH4t+cDHWZogrU3H32HaxqitfS2pzEEbTPHs/NQ2aO2azem1LUsxpwO
uD8M5y1I7m85v44W+Ac3x+DCy2Y7MQsXJd+p3QFQIOn4nAkFL/d2v3FgCak61ZBig369jyBpe0Lq
nwjXIjH9AOACc3zFyZ6PdS/miDIKi8EEoFcmTNXaWDQOQyCH7GuooQht+ebVrNehJFXLZu2Ml+Ti
9gO4NizauW+jTa96FGMjv76zjKjFlKd7GVhDTkA0PQnPrx0NbiLHGM1b0yVtNRiXhj9dWq9loaJ7
G9BCsBFCLS+2dHz/AaV+NlRvIyUj8JZU5s7HNmTSpSn1J4MaVSMy4Vfd8LmPDuJ1CMRy3/6Oy9eQ
1gxLjGBSGzQUjPuxBWkYo7VU5gYV3xp1XdzidnfinT4puksxLStSgSaOWSw4hjdw3vkDDSAbN5GV
kz3n273gxD4kKfGRyl/ugG3xNXV9O5kFK/QJcKBVRBckEsDamEMkJDWw1jw6WnP2htGDOs2d8gq9
4QH4Z7/iw/9kVYqi9RBKBvJzS1geXtQ4sutrRLQx8l22CEMUQnskLJtab+IewvIrF2181MVfw3KR
qampb1KbdIi/GWM9/UzoT0KnQ9ovuVJ0patKwWxczBhENq6cKmN9YL9H3LY6RD1dlXuqgyIDoenl
ZniRF8VQW3PoJ+BEAqCzgR5+mg8SSXTBE9wLyFVSYZLI631NesJtNURMShlFgoGrMjl5nsaBvxbk
gk1SDX6AHBExEyeH2ptbUwdnGedH+adK/Uq+kFcSxV18QzLh9zFLS75fSj5nhp4myZ6qkTNTuOTw
8T/pJjeKwVhK8krvShCNw976JWtRerBogjQ1Jht1j9hxCHS6rhvRKa+SvJsieqoI4911eZAeQK85
3nU+sQydFpn+TJHwNUJ9YeiQOT/07rgNDKLwlmK1alm6QwpDUUzzFm+eiJA3t0KMzkOdEwJkxsF4
GFxzaHzyN7xksApaxpVnea9qgA5eYClNvf9B4xNB8N5drMoNwxXmjNOyH1RQ5hA54bfPmY86XV59
UmYb0uiCrAEZiy3R5ewmdnbnoiwdGrWJ4QcuV/uHjDNgNuB6rc4zBb/xepaWjdAw0SLGd2Ii9bdX
ZIcUvNa15lwrZ/zsqbjbuzZFLxkBbP5wnsQYQHrwDAxBEkFZ8DOndwUNot7zX5DhYVpItM1BAbdf
H5+LFYMgjmMw4pIU3i23Ao5hQlMt90J4rOjvSJFyMp4RGK9jbBqGZLBOffCmQZJ9v2QNeneGza3h
ZtuFKsA/ePC7TvtGjYrU0BiCDWkD+2ZhwcM17NKNHKdzXkwRuFFrC7bfMmzSiWFOKnzVClZVQS35
OoBkKhTKr1ZIG8BPYc9Q6G2+OrTAdViZa/nZfXf9+RTWdNKVwohnuvkH5kjSq4OqALxBebIrnu1H
DOz7nZov6Fj4zUNSggyX+5u3ztlmVr0l5REu4KSew1NfzvuHDviV4N7PfJh8mK75tz/UQSRXpL/z
rouvLAG2Wo9vzXyFup4DbqkIHkqUqBKrdXc4OvWJl2kyx0U/h7s3ryTPW5Auxu8PoND5hO84wtgE
vJD9mx9t9WNcC8N8RvVK6ESwBaP2nWz6+MzWgEIfm7/Vd0lYmzCLC3aAKC4WQ+vYIVIot95S5qDt
8CnKfSI/5qW9OIkocPrFyUOnVIMzY30Nh0tjDqPORySdEor6UGf1koMCsWQatGBqJvO1MpsRt3KA
6HaLMdIU+9KH+yeTyJfJQZKeClRVGDwrrdCoVsZRxkXPX/qFP7UjfqDJ3+V/Q9MzxW8To8ePuoJD
2Roj9XXPxhYXNpTlU0P+xeuYWTz+fO5CdGscGnq84wJNxUeMsoNfIYtR6DdY2XR/CgRY46bFuvz7
QP5yTIfCYMTYp/0GUjmMUaVOHUKlp/RU+379mZuZa7WMVhkplL784+zXbx4vp74OikjJPrOzoHiP
T+r9+RfvAdbqkuwBJnUM2Drimd9EHhtrEjJeUsqplp3d/Z2xZvg9vtYMFT7beN75TRI6zghaGi17
skXfGyuTnuePp0077MqPjrZGsRBYnh4onC3Ma0osy+ANFxduqhYWpI4Vg9sK1M3mJtyB59j1H/ZX
MwtMwBsTKXB7gVTaP/0U8+1ys8OSA9atqLlYbO3XalMvPyFkMthOe6Q8+8l9zrGcbDuLC6XKWJCH
FQ6x7yJNYhRiPq0QvcuChAp+AVuBULGJNAWgkRffMEB1yeS6dhzBquN/fIMlgBHrao/Nf9YUaWwh
qdWY5vn01JhO2+5G6WoGlyFqkpjUjVFex8q1iGFioeGwDKXx0pLDXyti5WNOJq9j6a9BvXRjAdhb
2/Q2Niin+vomTlTnZKVsxvDguboVGsdK2qIT6ONulgjsh5PtmEd5/LTfEC+KjEfvPVk9fAqvl+iN
qUD0mqALcP9SteA5wHG+E/rOyfmB/wXhlqjklBBmbbOjwsSOvgQ2HP/T/Nzhsf0aWYMOfT3aiePQ
1zKmFfvgp96L8LhcYYop2wUGT+TkK0g2rf7pQlgyRRZ1gjUsOzNajaAFbTYUt/JkUh+NiVn4PzN9
BYtabagRnuzxDH34u0bIQMUUu5yp1tXbMHAOvLCwAsDIL8rYVUoagLuMM0wxBVSV1SnBW+7sUWjD
NmfCwQLI6HCR5R06yY235YhPJsm1rehsKNKri+lzaoHrFggIMb3jNnBxnGgMMpX096StHEhBsZpL
EaOCvCkdVIBatzJ/R9GnLWgoFrSPtCYCM2+74TLrwQGWhSguhUe74PFeoKD+Zk0XcJplw/cfqxle
LHjTrvPgzTmkzSdwZRK+C9oIvcWdLNubswByPECKuIor9ewqeOjnDKNLUlq46RCX9ejk+8qRz2K9
tcfi+5kBtC6tcD3bJm/ttESv5SVcYynQ8vEpkcHycbAbvQ5nPMhicWsM278rCf8uoj7YVRoWgoNl
6JuB637tFX8eFqBQY+FAKHyX6zLH0Iws66oIVkH9FpYlVgOxZyWx6YSEwY9j8sh+9RMCPqja5Rz7
RmcQEqiu5n+ujcq5qopKo65f+9BIY1d4IdX3ywexXHi2CeerfnEkTGDMrlHdwRAHzLxwGnSkMO5E
ATa7kq99/CO3XK03isxnTE2HAi38XiqxZJ6LxR6RCmy5G7ZjsvJrPW6ZyZgHeBgx60TEnlKfXUt/
uLudk8NPpd9Uy6yGyHn607zPg8pddqJ3H8y9loyrRhRbP4OKy0XJvHvCp811HwvqsdTvtSLSP/MC
1xq6gkznHUuv2/xQkUctIqdwj3e8kp8iPOLhvq+SAUDb4uKoLrr3rWBhj6E8AgZpKPmy+9GOcPdw
b7d2j7ONBuHxoDDtaIPSA7ETWZHA7KAmh3JCMQPY5ordmn56O47vFHdgok8kD950gWeQ8kcU+S7W
edatMuCCe6k2cp4wrWwqO6apIREfO6fWZYX4HGLhLhlzaO5xHs8Q5Soy4RaJ4ppTrmkQJGs7I4Sc
qz6vFBkanPsWYxfaqDv5Hvu3BrhkZUzDCVP31AsvlhmgTecSPVNsTF08V6zxXiYkVhAUZjauEyDs
qFdB+RaS1EWeGyvJn/j7XAtX/B9p9NMJijL5s+l83Mr/bojXsAgrUq/aVGXeSDBNBDbCfJbo7Jl5
HSF1MgOHy7QssCUYTBguwjIcS91O+0oNhir08bYlH0TcH66lsCxDLwdZsyyQJymP5uhNr5VQ7B5y
dYU/pQpyiLXLYqoB7mE8I3etgbk+nbnittsyiuvFHcd3tjp8a4JfoSWAdedcA9cvYPvpRPtaq8+H
w4ipIajvB8UJUHPNkYowWmz/zss/1p+MhT3pgfaHWQ4djcjN7EzHzSAKqL434imxTxKG9OnDMgLD
3oVJjA9dQlrv7kyZbSu1HIiRZluUHrDEvzePXblnMcVabmP+0QLeb7x5+cE2bsoHJ7rL5nwGmLgf
/kGYSN4iCWjbV2A/7AggY3hx0O0+bag8zsckBy83kqZN1wZx3HViu4Fh6SIF5/t+nwqCmbX4iMYO
pp7rxjNwB0BoipbCcttYeaFij9/yN/apSN8hapfqYPlO3Q5o8kE+q8+z7e+KfaKNcH6Xt6i+ldkZ
li1f7UfKuqCBVfhfiDBHMdRDklcAX0ASB1Fb3EfoiYio4vIhIrE7iVU/hhA4QHISCdmO5psniPk/
zgUCLWfbwUj0np5M2EUrXoh+xZHTYWUITJe7UJcGFM4XKltr+znL5FqOrwPc9o5Oc0fP5JVtnIf2
qdnfhqzu7D949Z7D9hB8vzxX7zB3Z+4ndBheiE4q/lBFQoY0FZ+AdOnZqXwuztKH20A3TCYu4Tgk
JEixzEXm7ZABSrL9PSJ3/08jPdEvOhHNG+SyC/TeRibJu0uGRnxdEM8v3BhB0+VBLgk5uJ5orxHp
RdjRX3X7S66XeGvzJHx3nBvgEewbEH00ixMVlWZm86rVRMbM1d2mpszhAx2yh/KNQoZwlT1afeQ7
bMy/nb+GugTjynfu8HtJIPNUHt6VBR+s4q1FBehjtigsIGlWDzy7h970UG/HKdo4kwL0D6CXPdxV
BsiaX6Q9CoozAmZU6I03gK8PzcJngNUa7bQKGsY4l8txgyL7Zwpd4/fkHav5fUuhSKZrGldQOcTv
plGSlu1qKEPiSC3y4jviamrxpElUTezyvwzvAgJDVI/p9abkYosb/rVZ/r8OZ2oUvVNV9RttyD4N
ihCTspfU3cTLYI9wh5T3/7AMr0YjQRKyvcNDZ9qYICefNPIqAuEEb3aZBCfZeYG/zrSyXd0n1eH0
hmiIjZSsndx1dUmyDDpE7OlGxHxHifq1lf2IwOIm0TdtYr076ptb8STGs8qRDXlOIpVnJ8hF4mm2
JVQDVVrBNVJAgzAm4BS5HQ6jnciZ7DZuVof+AK4cuPTU6wVmM+Nj34jzTq32uI+tbowaxUAS1HhE
PN9dgVHeuv053f1LqWB208TWEm/bBynxoyBpsOWGX5j0Xaqv6fFfEtfCNdq3JqFhVkyjOb7sJdIc
Tp0e+SjdQ34ZvfSgEUzEZGGfEDlqfgk8JFxqwYDwiXOCCCV4jpxRDoUacZzTGjTTSJVcMD/01bL8
6WqUOTKP9Szut7QaljL4X+bomXEJfQRTBt9m4VgBuGfeJpjrAldWZBKOW6+Wuk73sxLL4RD5TKaj
gAvkZ8eS3rH6zrJ7ILND6SNKY+i/t+lMiKMqmJl6B4nOFcpKZM8en6AHERZjcrK8JRCaZeMzP5Hz
jI0ymnRXidlwviyQbelwqiguFYRXw75UtzHzGVo8xk1t3khgMsUFrhxnzEnTPGrNEqatwaUhPgM0
9guQHoZR+JI1hC0rgdLdH04h0fn2fIhAc3QLcPFNAIIfIg83A/yuoHJIl417TgpXLsGlSLp8EM2h
Y8IEHnVg9HRweijHvcn6PRGM62yj376Na//JUtTM3QRupEVBHferXK/qx/ZXbM3DHMUXLvU1ZzGV
3fgTmHPMIzezJRwr6us59eCs9Bg1bsmmNPn7Z1yt5MnLFty+l8KFblQEy3EuL6U0BH+pzxJLm4lu
UC9D5Hk9BLOnzDOmKGe8sUuF76n5LyI27XGP5L+0DE7l5HKYBd5lBCiuTvyRSrpq1M1556hrURly
gdbN0vAVvQs/e4QTzRvHYmj8TyeKacsb3FBZZe7sr+1orvfvigrW6Y1/T7aR8drAqIsdG9ellfLk
UPhnnDg3WAAa3hLwyZBJ3dG7ulmnEc1jcPHtlLq7sdwpE5s54TVk2BcIN5NOVJuK6icQJ40JSO3P
t2vcU2+N09ofYR4Agw57eECox6/KRDCCNtjsUTm66XpShOvBM2tVq+8QsLjS5eP46597+RXt2Yo0
OPMW6qyIWxOWg2aeV1IV+1J5x5xiWQm+XVLh2+OfT2+0cN2U0/XLkdimU1RKioHo+L1Rc4VSVaFR
nwBKQXWdRqC42k1ize+3C0HFdVrKOhZK/NVU+4qU1+dh1spiYRjI313WpFr0V43aqx2h0OdRMMH7
iJ7TtPY7cgZ52PsquRzRNhG+kxrx7mazV8BLYYNYABDidSo+Lb82KrHAMcOmkJuz9T71JwkSiqlv
bWoAA4rnK0HjPBWOe0kK/CH/gYOG5nvESyhg+6Kl3AGBFlY06G1XuQlF4Udove1GHO4830GKzg/J
b3+QZFkYZqxZak8t1iKdGRd3JkgQvKg7gNnLF7a6W/6bvz7eRhl/jb9x0mmd0qQbhWbbvliB7vuw
xc4ukROdmHFIFgpMu8f36wGZ0FsT1BX9nBsok60jkJzZo1wYToHWWhVu2pNk3jEANiq7NQ+pRsx7
PCiSzt16HsxuyFkZHzIm9C8KgwFJSgyqlhDkBb1fJbujwmt5/wr29rR6Mt6327kpvD2bD7NqVs2T
vNLEly8w7tzLZFRjTC15LIsl4JF/0oacjO9pGSMwGNXMTdIUWMVl/ue7ZT70L797vML8psH30k6H
oxmewg4FkxLszhj0pcGjmyOZTOGC1I6GWaeAUKll5AjChi8rXFZN3TUU7ebdxQ72/pAnqq88Y9ci
U/HUjoX7H0QSd8fV/hIqOeDLxO6eRndo8VeCV5Q7Sp/9E/m2XWIdaDn6CKg7wjQgGB3nzsrFCBHZ
OstxREk88dNXJbQvqStkxWBXD7mmBx6LTM0LXGUGz1nXVCteBaGcFcC1WkyvBq8K2S7DgihkPnEo
REYeohlI34gWHVkNthQC+W50g2kzhD1D2h20tKi6anBKwdLjrHPv0kU2ClPz2/i1Ov//fQFlz/aY
gQaJwDMbFrVYV18sT6RmyS0fjaMETN0/PCB0fYSYICFzK0BjNltSThxLudTZXTfTvsOvJzUfkBoL
2tewSbkulwz/Dk7qvdBB+brGYSOmema/dcoWlv65bc2P6kwIKh6BYSPbUj/uB9OPLko0XzJpD9/N
7TjNNyOu48VDDsyDemfyaroAXVHejkPdCgs9gsbVuNG9XJ9xWb8vqtEkT9SBTvy3OMJB82nVkkPT
aM9M2etzCapFOgHq92ZWii0jVn0nl5rFh49xlDLKWzHfH7Umh0a8OBWFuAWmf/UxshMkU4auUBIc
RHaOy/hwhxCW9WGVvVkvBQdPlHmMjfaICC5efLIPhJg1Yb+zv9+kku9QKuyaaMGIqKwYXwXiMYm8
Q6qfMhM4zYRubgs4gGIlxt5vHGj0NuOrjpiaSKp1HrujViKEwnSmErWOIRSR5siMrgDz1M7a3mJt
HCWQ5GPSakibuiYl74gH658Bx1du+wnddWAFzs5A43BDLRlJ48VGmqB4dFEYbf/BNijYwq5fH9w7
3eIJegyE3aea78B7yG4XIskXN26NFowli1X8iR3q1U55Qz8CwCGeoYntNm2Ev+WuissIOuDLlX6C
zg0K6hRrOaNPewjLMMIcdSNRXytiqDyzgGgfZSz1pclotNMuVVsjMw8mpsSAihVdwIPSUc5Q9nTd
8cKnqq9WvsRj+pVVhdtp1GCubI4aXODRhjnIDRkFaBRD2OxXRy7/FP2Y0TPVnDAI1iaB428UdT0D
Yg3/LRcqnv7VxknfhPt5yPHCvQYVk+9TcXc5y2b2vEIzpXu7nEqbq1mejY2cih4/+YJfoVGhIB/Z
1Qe7F+DOAUMEebbmRxqfjgBK6LpWVmADaw4zrTyRTl7Tw/DKlWksNGcaP2844v/uk2X0aorP4jFd
yIUVsDwT41OKlk8fPWoD7GbgBC/O034pyZJGqBCAsAvqaRjgvAx6oOCjdR7pwORZFzGgo6IrlEgI
2ElH2WlyHJCWM8ihscvQrKPSvwj04J9DcJhX4N0WN/P815Pnv/j/oOTIs9l5IDnBCHdTUqsfomep
RzrtWf93TUnEckj/yXS0iXCqk2LXNipXstI7PwdCNxVQwKvT/PT5pbeeyiXchssDTN3I3MrFAEmT
WIVGHhihtObKUvUGBEVdHndvC+7nE9G0GGkCxWfVcBw19n7R0g7B3CbOtzCeKcWPPXHbG7F6KzqW
iNR4bww5itfPERUAtqX1PuJp2NX7g3m2z9NOcemBYmcOxTNIYzPItANr4aW2sZ6C8EMma8sPCJvv
59A2at/rH1CQgyH3SymEOWLbgT/l6bAcuiJ3RaDBQLM6DsIdXUgy7ILxXyVBfgljYCXklOkLmvN/
V0xYqzw0TSQRT6XtaYwQG4xX3vPrUwiuKJGmYldZNeM4Tuy0cH3Q/ZyILeCqVq1CPwrmtWFRv0IM
rdxanwi6Tw67AAqqJBbFb8zvxJ0OXfHxEdT630kNxY3qeGXwcy4CDKwT7WJj8hhiLk+aXYJ/2cE5
k4MH8Frob5TPSE5WPGbuVupX6IaCE8KZAhzfD1XP3rb9o5atArYPbEeEujfxD4h1Ax6AvsRC3ez2
8Yh3brBlxMeWtqqi23eezjzvEtyvZU7THdaJbHt81G/XV/QIz9AkvfFY65+Zr8GWlvT+hE6ew94p
nnosZEWdCYiJ1X2TTlGHW7WaHIG5DKlw4MR4qwIP5Nog/meeEQXNoqetPgTkAHN4s2O8RiWIV3Or
vK6kRMekndo5eKo/6XquOahVSFlx/iG2ebXarxKxcHXRUSVfWtnsp8UOaDnHLV1pgHTKtGSMJ3op
kOhO9jlx1lV36p8KkPGLRr8SRRiBNzYD4SAjPIU391KcQEks6J6ibREbvFy3X+GuryIION6nPxP4
K0LPdMFdRs6iVX5cTtdQxIImQKCRIWlS1pPJv5spD0yXd44KXNGuaE/D2VpjpNr+qY9v0KcKL9dd
ncIzbRGDdVGX2nNDJScVJQYnW6daAcntlYiKpLH0IxKogvwxJ8ase2ZUyblA0wcaS7gf4+NSDwTI
KnAAkfmm7qPXM4I2kBV3qE/10aQQPVLwv/0s1NMbQ6TmCw5J3FEkVBNBkcoiyiKOwnoylMe7WVth
fL09le7FwvnOiF8auyrsj/g3rsOinhcjm6vixJwmwDs/K5bpI+d+47qNroz2na8LY8nCUzEIc4eT
gy4ssBTcUuljkJ0QydICDoKM0Sh+rHM1TqUf85TYOtm34whmE6gKMtbz7XJYsMq5sqv85imVpab6
ml2nJHbBobBtK5sIYRoDE+3At9PVHQE8F7yBGJuJ5II8VSOr107I1YYRq+pi/4sqhksLfHD6Re/U
IPAgnPr/+XtBq5gq657j9wTGtsl1nc/vtF9KSz9GdaMm52JhpaoTZcqbb+g+pAeZGq3cCUz+c3mA
tQocenP89PH2zo5GDwfxNjqUSn4gtWenM9k45N6iEmQLELBpl3Or12OKHF/ChE3KxioMu1WWtYo7
Vgp1+tnEvjg12XoBEFxeEOhvXLMq/he9J0tN4yvB2Yvbs4C+CctLFhqVQasbFGcUsDdY6SFbHxCJ
QkJmu6J2sLTnnBc4Vg/AksuldLhJxsHUClhe1rVy3M3WbrOiY8oB9QcENeRHajG1uL9hRsA2TYQ1
JdOi2QQaknOSg4Hxz0Jd8EsBw1t5lJhDryCRz9cOZUwc4c/SYebXRYX8GgZ04IMz6X5hr0QYln8p
e3njW4xbok66feYPd6DYA1aMGmHOFNQb7j+d9R6s1bFVJDeImcfK42E1ZYb0MZ6DCPmXejrTFHE1
LA6Ygpv+D4pKOT2MLj9SkYYaLnk5ZNt06tdGZS2CKef/m2SVXOf+ySw9vWCtG2nL/ObGi+B3q+WU
uu8FKYfTaStFy9/rIGzkxKuarC9fx6XdYdeRaFpD/oeUeZnCHHxrCCecbELhTAqG1u5hnbPIXDab
lGQEiL3dWvzFnoXP8VE8kjHRrC+XYIT+hfwuyZU2XcZd3C5osKq0h18BKHAC9KBnd6WXPRft7MWW
EJTJwNui/ITIKO+KuGv8xOfaW2sq99nH8I/tdCCHkU6pA9Ua41jHMhuG1E45KswYaM9MG3SVTAN4
zbDAkfGK2tqCShIM0TRd71k5WqoUZVF0tJJNJE+32jwf30ax0yYlUALs25CC1F/Kc9nuB1hxulTf
ZPA3Q+S+w3h9T8LLHDdXgWkA5EyZCmfZfSj5BQbnn8IwEMn4MVjCQF81dvY/oaVbhqkRMnnoppfU
l2W8gQTg64k1DBz77KhQfgWk54YIEr+mGnwXCbsj/2Ll/+pDFsuFd4peaqR8/6J9HGGNcF4ZT1rh
HPZuAcKIUnH9bKmX1OpNZ4j1hi2zbebQPn8ljOjHoRDdQ9njFypx/3InQuVbSlZqQIaKfZkWXORY
yriTLPotlTfJ+aXMClo+aaRg8B3O0H4u0i5DjZ5aIavjnhRjzZUayBkkjIO+MkI6O4ocNiib/C7p
FcHa9FC2kp4XwdslPvwNHRK0OhrAfD3/Fo2/pLH29FArkZ2PIow1xgqqY6AI96OtbeipXs6WpOds
MAVO6iG+zAkQSadjpLjJ0Iez7DALjZwH1DNMIT1/mGhqF1DER6NDh0Gxkb2hc8hPzeerax0MRCDn
x9UwJmUcAtM7oMy7ZMrEBCioKFDaLmQZqV9PKhNW22InJkYqOVGENzne7CR5jtjvNx3elp0qPyPo
9UaVZucHt4y0mO/qjdSdDVb832XpXD7vD+AxTjHJ751iD1ph05s2uZ6xVVBrxHCDO8rA0zm/M4Js
D2Kx5v12gi84aaboOeqwzgsz2w08xiWJE9Uub5JAE6ow/WQlemUelDf4z/750P7ZLxL+8Vy3xVhW
1O8hrlsqIqYkESU/4IS9pW/A0fXFuUUajDBhNu7y2ixN8IDUvjJ3Q4f03ISy/eHONDZCCBBjAJ3H
O6VB0wMNFW+6EZ0S/VcELe4HPvxWZxZPuHDyNQB7H4ZrMDnTxEjTCCeF0a6jo0TqR3kZ/RrPgWD8
D9Lx/Pksh8PhW5GEieNMqVm0TiGi4G1EgWks4F9D5WniyHdir600w05y95YnjeHanBEusrgT4ERM
dKMCk/uvGSGZ2rMUVvJnMkGNWXkRlRlQObzZmwkyt/A9Z4gzUZN2WFQNmYR9J95faqKWVfLJkaLX
LjQ9MZVYhRey/+yyCYlNC2bPUO9TKm9aOZIW8d6uWzM9V0xBHerqKCM727CJNZ4DshdufZP/Q3jw
zaihKkXaWYT5H2UOaAXWCnk7yf21eBv7xqEn31nlf4CnLkIU1GO6Zum/MzS40fokL7VovntBVev2
CSHdmOSHeeu+r0NE78nIyXSRIHj0C4po485pJ3ZCZ+1OiSrlDil05S77ZbMzuJQRf3vDZYWGWfx7
m9mIqBG0q2+Euv8RstbIdjFVMM5RddeI+M2HhYH52uiZrpLL1ChbayTUgMbHUOm9nSKPAeWXV0+q
kx0BA3/RLV71Xxzp1FCWBeJ9haWdW9y3Hts6/qfXKc2KTrkfCaL7IKPU6MVhcR8i3lXW224LmeYZ
Ueu0DKSKZF4W5rf2G41nL9HJxc3XahXPYJI5LJiXYWHCrkZWoSywrpGaFIfanEIVFUwKjyCoMumj
DXmdA6ica87D2WLnABhBl2nwyKrp8w8rCombzzQFosT4MmnL3M4cJx36G98rvPBrzinbt5x50zPW
nhqz2KDD4VvSzD88RxGIso3xqhuQSVXmxPhydCVrQ9wM6RC/kH1L1Lg8IQtw+58BfHm+bNvQdxL3
qyvUaQR6SrOX1At1jB+EdTIplxyKea8EU94uN3267NMvhnKGT/yApxwnCga5aPDYe4ZkSJCVSZSd
Xk+zukvHqfE0LAR9hMxM3kzFDHay69eNduApHSIiSQjBl2dcCppO4lxQVF+r8KPrLJcQzhTD6SKK
BS+uFJiyBoqbOZK8ITaTos2xWfqfK237FZKhM1zfHPeTXfoIrsXZBjsAZsQ6nCCM8lS3Yl1eBtZF
54aaKef3MEMeBfwKQRA4vgRj+DxfvLrpjTVwVm3ghoMxSa7bSEP5g2aec6iKKYp+OSs+R9mPpYmH
XFEawLCK2rnBJ9+l3DYAzi2YD1Q4t7XMaO/yOkJ8Z9gruNsPybTIpYhZ8ij8m12uzR6ODdg13mp+
323s1FJb7sdMTDRDEpeaS4rSp/FC9xs/IuA9AOvWY01IilaOrCqX5Vu5hc3Y+8P3YY/0hQmpmcct
eTJXyNqXt0Y4TCMWAnC/gaAgk6TUtm6jQGEci7MDmjbBFSvp4ehOZED6wQ9QphfJhvOE8ylPh4AK
jxoGYQbWK/eQyrAMHSgpEnQdPu71rVcZqque0qOOKCySodr9YX/QvC7JpCdL8LJPw1E9TDgFz0cl
AWoMMrawAPNx+hi11NCY3R1IwNAs5j21dnGrIixbQqjNdOqkgMXKJ2jstMHWld2L5DMplAU6QKtf
M8A3fGkZ9A6haACK0B4Vd28KZOJ2fqBHqWqa2NiUJbHbwbJ7CiyfpCDZKM2KPYhViRbJWry9wSzL
8lG9IQHuIPI3TFR0VnonVC62KvOzTAiHLyzDAywUHSKvUTDR7xaNoy4kQVgj0Sa4Fv4r5DUnNgeX
nenlv6S5pY2ZO3dnBekS6B92E0qU7JowfMF5cOjLKTfljlUWoZLx6vLx6zPjuzNrngJBhIZLCVbl
5WLtf9UD7jzf+fPBq8lCwi6zf19av4Z3zodFS7Dq8IKrMhstGzB1LbtH/9eOI3nhkZxKVKCbDbq0
WTa++OsYEi0ElrMBD8raKkC2aC3qSPEK1Esywb1YmBt5XIuOSqORQ3jOQFwhOPHOYz7njDvI0dfW
WHa2KipW0n2AAM2blxLAfisxy+on6VELhKNwog31sJmzRaTK5DfPs1buDlj1vmulgQPQ7U+HuBJE
ijqoE45kkyh+2sca7DVOxQTnA5Ii3B5k+5hTpxiAyH6UF/LHM/Gd6Y/Yetx8CJUh2z03B82sfvBN
vYbTSwutsL5bMrihoMgwJmMzmEFhfdcU4F6whZ3wXK+VWs4WSUroAC/TaFDHjDAl+CT1euC4B4QI
tEq1yjOZTS/rTsKuUNor3KyEWumGyc4Wh/nIJXT+Mz5kIsQFDoOHf3b4pEIsBCvbC8NIxtA0N4nJ
ygvGyz1DxDXSzk0/wmd/TSJTvsK2dW914oJ3je0b9G1XQJEacbpaVXEeHc32Lix4PHvzz0zPVJVy
WKnJam18PYFfmsfb44OPSgcKrErifXN2XxoKMkdMaMJZM/XDwFawTuY5ffoZmD1tqO1hlwSxN190
hDSvuhRaZlLMen8y5B+/bXm/0ckm3P6mMj5xjoFKjK4lHlCo2xiHZ57cNhDwTbv9NxzIA7Yat6Kk
j1FJo0gAigpNHvfFbyaX55IKPM3IN7GEu/5Y+8Nb8UUj8W5HNQjd5KLjONnGFc7RtmHoMZpQHbcz
FXwbz/njfDtY41IJ4eC7OihRKDuYHGLVCjweM00GuZborbhybtwJAr+Z24cMKlXyd/bgvhd3hvOi
h2CpCb5GPcPfAt0ZCmsLCB+zvLZTxpv1etQCq+VqPk+QtziSPRV+uXJBb5qhr225TLDqLOhGgTLq
vxMlnw3QT4+5V2Te2yuiRHJAs7O+jzFt6ML/uIiQMrjFqO9AZcGqqXj6701CTNlZIOpGnKWjT8ix
m8aNd9XzsCENPvgnl0ETwPl22G9o3nJcHFGuhdu0CS8ZVAs4XhTUnH9F5gTBmIFMfDtcEdRBKQLR
xnOad7EJfX0p6oRGdJU6AVqbl7ZRbINfnNIzs2as2CJEFH0FVG1UI9Wm49a4zxzAqtQO763hygme
hD526r1zknxXxFFCLGR0exrK35580/R8VAR6cxXYt/HN4RTrTAVyUQIKiSWT1G+2sU9Vv1pRDPd3
xnVqPAMnk9jnIEAI38ghnMizGOASorqSCHAOyKVFt/9cX8lmlNZUOBWFwPtEfXqlh6eI9t8SMdL3
A0ErsG8pssWDCJ1YpLwbd1YNHdqNzFhJOPUVSZj87QfaD5Po4iKgiT0i9rXdBoeHY+Ss7gKLnzsl
6sXl3DFlLx0bXnZW9FDadaZwnqNLukihUlKgCA84r16c4DDSlh4+iyko81jdhcOHfYMBbtWAhdbl
2PGPIOxj6VJ9ajxoLWWkCQgXazHsRKlTvL0Q7fbypR7eZDHoO8+oDxe5s+9pAqe2c8DKfJpxbHCM
rgO2sXpm2PDcg9GWR+K6jdvwFNvty0FAzblsg2w3VVDiNIXxZNpQyXHIz7GfeXt32e+3xCGfBymr
D3hlTbxSmAJfet2QDpWt/H9dRYhseTH0hKnvIZywCOob+vGgMR7RALRvwu2fDYbnNapV0qnx5Lg4
SOGg1LmNpCLaJw8t/7rP7Rr1dyJHmpomPcktIBJ01sp6roxQjXwKUfyW8kJHsqixKXoJXEHjV7qr
aEWJhmjx7o3cXcKuJmWmz2qFQpEhxa2tlfIcpwwcaL/D1uHKM4xSyYO1233/crpYPle3hkRqi03f
SgbuDkKLE++DyY8UTA7AhPrvwNLNRCzEPs6I+FhDDIBy0Znvgywmke1H4YI6Sa9DJxRmuDBO9Gty
irOPCIrUL2cH/r8v6VJf/7TiG3/TUKvJM+HPZAkBbWJILdlDtnM4mh3nUjzriNkOitvAaCAAqobm
WEnKFes4cpS+PiKS0HCfyrxweGRX7ohNM+xwnjOKX31CpwsmSEOlykEvNaRgLORWnWdGtFZw/FDn
2Wa7hILCHmd1rl3RBZx6UBOUe3xDPJSNJogadCsz1AYVo8VxrNlvJTK/NZuyONwEsU0jHTacX/9Y
rpKXRHPY6ohIBGWphOjN7Kno5dRwDcxybcvpFue/i+ivONN3hp8+HnpKdN7uaH0WArwqkT7KVspA
B2Uml3vc7mVAl+wgVIwXcmBfA4zPAbSKo65Z3aFoUL/7LEBrSYUteWe2Sz2PdmXWwhT/W1vyAsWO
1S7XOsETh7gDCaPaCzJd9QhRAudm5J42/HxeXJf29uXK9W5iYGXqIW1yj2EdL3YEXWl6di+SBclj
RUVPbsVcOFuAK0hNEGevCPiu9dZc0j46+gHm3n4G5UkzgoABD6Pq0wrT20KEI6HyQQQ0cEwuHddL
PigbgQ63GBvpXyHajqF7z1j74mI6l45pNlg5JqMVPwZP2/pTV9bEG4fuoZJn7W9wr1XTNGR0uxyj
4wvbkuXZaryWR87tPEm30s/PlsqpYTgzP6np61JoIbbDn4ocm8Sp263HVqRLM/mesWN7YnC0Jhyg
kv9DExGheijUk9TdnIrsM9tJDT4XqrazFzNA3d+OVKcNbf40ETmhKivyjcvAobm7TmON1ciTY5ae
C0IEiNHZ5P3/EtogsYBmftHPquDfVY+YzzWXoUmtdw1CjFCo6/mzusdZnq9Fv7fCZJfNk3RPXlYo
oSWKjPHcRdVIfS9viciL7+LGgBzcO3XzWtViZJ1kZolLC9FNH+rY1bZ17D8dOXETNjiCcNrio33w
Wh+Ybr1pyFppazmDVC7x9Oo/uj0lVHSZHzMMeV+T1dc0OBusi07xSg20P6LwGX4K43TAQvKP+b5+
Tmyz/1AoBTwTswhuNPh6XIq84iChhueaY5NdwXvQcPmv7zjFZWFOrnEQDpx04OLvyvfpNGqaUtnD
1xVlJvyKtAS15F4cFGfPwEW659bqCLcNdEsLeOsbwGSC3lA1s/KzERRU6iqG9DGTfL13vKd5SKfP
4pAblZuu7KH6nZRmmLtz3Sbcb0rrZ9VC3hGj9IEyKD4j1q8kq8xyh90vJ1G0Pi03jEDFZHOW9lRV
g2k/Fm9KVLusrCaSGUD51HstApXoaBqbyHfN0nMjAfXo1o669WaiHottWvTMH8408pXWWWLIppAv
M+w9goU6PcBJfc22/C3gdzoD2/0+ZG4bcL/2b6LvmeHbVCsxfyOTuJADu/en116H5BKAjqKjFRYH
DJ2tTIkO/KrrjNBIzC1Ut++7ofXnPC4n3MZu49Ddt2Z1jSIn1j6KKN1iYQ1GrW+ZY4SYI06y1smo
2GAiGFQ3EgcP/Pr3OazAQmJr6DRffUhPeQ/JznsFAW1VWSXxYuxgNLSpmCxVevHOpFrHOro4CA7d
BIZixJcKB//FcwKKvmiBczNjrfdTzxv91mFdt/qYPNAzCt4Fh3jZRaajqWUBTxBvq+WsAJH7RfCc
ucsK3nwp2tjJRIOPQD2bb8+Mp8VycZI52R2OE1b5fGkrKbSPzvzV/dPCH1weLNNw3zh27DEXfUr7
m9TJSjvduOSxcKJ9AowYiW19sQnEL9OTVkcq7d499Ac24rJ3cQaogxUdQVb55OuTLtZO8BNgGkCj
X9HZzSGwv353EjIgEvMAtbgwebXfQK5wyVpl72gjqIW8Ey5gsNP+H05zkeIFcvrgVhWmmwueSe9S
zL9RZezPwQ8MwzGSX87dUwdjA6KNu3uCITCcFS/gYeKJf8OYsDzsmJ05AR0sQ90YDGLK+b+uG4FA
4S01/kpJNp+yw8I0lAGFCPGlAxNv4r2RENth70fCkX6PV8IYPwZ7b+NzPa27YKDNbO5XWpYd/hwl
QNgCvLgG5UbFKoWeuTyBEc741xUEjhGl9kzMnb29ZWUjHyaKMFJDRoOpZ8AJ/TJO/n2KG0XsjuKt
HxmoudsIymkVIptwIILfRzIx0+3RdGhLc/xghl9rrqqv7EsEPDravLjd4Pyy7oUZcAOaFxpvKSe3
xsJxB4DaNXnADgV5pkZys5/9RuhZcAzc4iNiQcLWfQ+5m+dZEHqRfmO0tZRaLY9BGsnhaLahnr5D
5PnJIJobZSjX8Z/6rBF0bw0emKJhmGlq2MiHoOS6xCT92zCdj1KhUc2W+NuJF4FuXdf0bAb9nfgE
+rKVlKV4MEyEVmLjK/MYC42T3PrGbPzUKw+OXTnA792ab+3UpwfKewhziPLkVXhvcJ3mP90QR3G0
+brLMMxUwHD+Edzgb2eMqSLrpydI4KKQ+ipPnhiWPYs5YVUjkoO1Z+0uRIRrwHmnQEbjN7gMo4nY
luxlpqTQYTQPmkpFOFOjmKlMAOuZywfibMaAiZTLb1OEMon1+9/Z+IPy+fuWUFFL3U1tTKrqUwhP
Poj4/xf2SGAt6PJlQfDPcvApRmmfqIwIecIyrOruj2eap1wnHBpkJXUI0IfhTM1Fm+I/X2LhAAXo
aK4jTnfaWZXxH+fYbJXazHIGUrr/dcKVpJgu7KjhIw5sTDPI6NMqSAE0Ns1KQYoKsazy18XEn8F0
mCKyUejlVM7YYtXlTZvVqVcZKzJ4dwCvqYa8R0McSiWUP9mnLsdgFdSdFJfpnuMrlDRYi0szTajc
azUST2FBaQy6OQd0UvEu4W2/HXer57muitT0lzYiESJ62jpalVz25kD89CGw7sI4vT+EaYSrv+Br
q+dzkgpDD6xwaBX9uOGc3dkBgvm9oYtNeUi8JYS2h8GY4WU9r0h0oZjLrVjcoyqsCclWWYGYFw3o
NEj3FEM5edbVdBj8heXhF5Y5WomW8ukt1h0cEncIK3B0yDONCirdkMPv6QLQA1PnEoiXVVo7+EgR
9/v+shCIgsYPEUByLuaKqqjjQKA/dkz4ssTpe/IyV0souHXIxuv3a3PBNeLcQyajknMkrHgBKVBD
dbsMcYqBLTQePL+stThohIj0tm8iBFyg+W5XJITg9NixbJKGBb+ECu1eMAAXhHzzsTp/+WR5U65a
CoAFl282O1X1IK1jeMAPWyoB5K/6LUZrFNjA67wYfU+krhupVpmCig02D959aIcMMHuPXF96LDGq
Sz6R2WZGJB2K9QTBC139FVo/QP122qYxpeZmfzL7r+Mn7wFCRsgqEdnTd7cmbW8lLRY5qkU7yQqU
zcylkrIVAJs7IgaA6Qbds7StCfcRBBXbAwPYdRUlNwaGVl5Z/FxUYCc6H5vG542qAsiE8oH9k2d+
8D2GnvVcPwbGzM3tBODt1vmJ/av6KJO+l05lms7Do9dOZg6ZDFvwfWuGqmlNG8L4hDYT2gaPQ0sZ
FHOLDojzCNAR0dw3SCgyn2nb8drXAqBNyXo+DcouWL6YRHnbJmR0QKV57FeSN5JLRUCTULinkuXD
4P4nWNhXDTtifWT0+7qk9pqNjTf38kVJOwTCZkurgd+rpKFDsshZqsSZ1yAgnYloKt6HVfA8JRuZ
HMMgCC2FVS45xxGPfKtH5kb/az0s+adQ36JAw520EJ+XQHn3b4c/YM87K/Sjw/NgatBbM7ALPrhb
o9fAVdmGVyByToD03CZYXseWhF+U2l2rKd2kf58ETS3ZojyLPAiXU/hLrxgA87WTwpr7um1G9m4/
DX58aRFtPOS58uCEpwQ1gBWj+p5fdrgKytakG9gVVBqXNUx7jtr8/fdAT9VhJFkCUCNqDtaIEHZ7
h0gH4ESqABu5/SqcebcZrOht8NAhb6PNlh03rFYA9/h5U/gLCpazr4S8cLA/u24k7u+KPIXKpNC5
/mixJrMqMWPlXrEV2aydo6LKig4d0TP/7nxltgNMBF2YnRrTc0KW53ucOkZxx1L+k/Z7kd/h1HsR
7wNnvPWPswahpALAzIQkC2kPp1q6n3PZ4rPfK5RtrWRgmTcujS/7BP6V29g7mI1bk6XovzxOtEFq
MLxK/EVYX5znOxlcgPSU6Cu6XGTV1B9bq9RYrxk+sQftCs6dHKL9k1PMwxrdIPR6ed7YS816XYin
JI7LN7Mg1FScnyz2ZS2dzQwqFL6/grVw9o8RrYprg+WKkugXOQhYBsqdEjERL9Q36pqns0Omit7d
HBRXGPldbLL1ZVmpzyT+W33TL7GbqeZsx42Wd1ANt9PbJ/jajLhPoZKRwsTKh+GdPDgIibNg4VxY
70hNAVOvk2MJkfW8swXVEgrKVsIGuIix34gDCbWaNkzKAtSX/w0QQwfIRwG4Krcw4NzP3Ancqczu
b9KwchbUjMC+mKs7/uJK5BHBXCrTWbNuTT0si7le37PzbZOFRY1p7t7GKksNbIrF5APIHd+MoMli
M7PC7jyTo6E1w8qKu/DcPgI4xtH4vJE0StcjsFJw7ZOHI4T6Vj2w3yeiJEblXCBWjMvbXTBY+ds6
/6yfW6lkzJMmHJE6f3WlvHQEd9oYR9u96n6r9xR7EBoR7Zu3Taj6mHSRw1rDUFnF97J7PKRkl7jk
QADOSug3hrrSEo20f/WY262Z8kXj/K9hcFGrWf4FoR3fw4OS/JsHg4OVIceoUy7mYO9ZbZZBz0hD
8/b8aT5v1NOygsxgyplpYAxvgeY0ZfmUZy5EgG/cBlJuBZA7SLVOAsz0YIpJnW0fbRVeBmims/UV
rQ/IofDzMS4PGXk6wx/xdjUZOAAC+DUcMtzt4w0WDc+RLp3ho12X7JOEsSHeImYmH35rrSNxnphC
H6oLhMLGeb4sMWSR5+kkrkpcfFCE8vN0np+AW+FQKGq28QK9dK7mox+WM/IDoghpkKp4GxJFDAU2
5DpqXlErW0Q4PJqsZPYVPSAjKtoeBN4DwDScWIoZztX1qWZrOTXA3Urn2xTgq12QdUwlOFZjO98G
aI0AQfxOcPK0tEO8/cuB4dnYU3CMLvO2FSl6IwMLNYUagZNZpRgFcsvEpqGAYYiawrjozzSIu/dW
Emv6XzSPZ2mJv07dtVtoIMYN/jDxSDnuST03LioG9++kFjYljkCYu72KxADKJrckdn1LE4p78Bva
HiRuxcPlCeE/Wz3KPkNDoilkZLN9SU9ucBKkLX/k69xyYS0KXrijyw9lXy6xuozjCqbmQBBlenPg
um8y8s0eZAT1qDgRLGM9adIni7omrKTeEmvOHunCcoFKfdJLv6CFrb8TEEfcCBL+lQhPI94XKgn5
IRpgkXiWUcWXC6qtNVPk0bkpEm+XgJwHci1Si7wDHUBse+fKj1QVP8yqJsxt1TjC7UZzhWZG7jhY
gcy8eO3Vc7RP4vl5mIpYUZTPPm3w7iV5trlcXVae6TxEnMWJNRNIOQLH9UO58+z31rXX59XpZ/NC
hbV/UsC4+8UQXgX1ANHpw3uoBTAEmKMkyCtfa5dNDSLzUKeYfLtpxYlrEOX2IjWnLiSSIzzkPQ+W
461OWoAt7x5WfRzlW7+OrTl+7fLIink6gyZdPcStHQ9JWjysvc+FVhh0K/UTL42t8FUECBWqS2fE
cmMhJuyIpigTnlYfdy7sRcFqEA0qyD0H/3ppqdT9jK6rj7SohAf1MP8xlSYHJ7nEtDlbhZaJ+HjB
UyOmfre+zKiBV7Jjg2l9LZG6uxOy0GQWq4LMfeHHnetvXyYW95Kqc+Ikec6CDguvGqHBhu7vp7pA
OD0F3xVN95vG39SoEUsDBLDFhxlbFkPZjfIjaHSpxgRHNWutKGRgXsUXXbjO/mEHa2vSVHS1ZEIZ
Wv9Tf3b02pRu5a6DomYcKvq3cgPr55Eu43kPLeiiGOQZNJ54mjizK8ayOpE0WvN+3RUToyOanmyv
Gy7GyLRqCpzq8yZaUcuabM9RB/rm9w6edRT02ekSEUB1n4eU5IQbNjPfjE9lx/SbiCihx4AHAm01
wsFwYM0onYUA2UaL8WwA+osw970zs75pvSGqtyGdUPCw2TVLoDaFw77BIkT8P3wbVN+rCDoGDL1F
p7VPLDenJEQLuu75kjCkMszNw+v5imMx7UIKH04mKQ6IAwI4ccTTQrSi/CMV3NotmkocYk5Bltfh
n99LJf+JejD4mrs+be4MpsmwVbsPS/LzWDJUbfuPdjMPXIucPXnbU5AKd/jQ8khTAOk0RpuJL3uD
S2bwd7Kc6RyLSB3zYq04ASaSEs/TncyOrK4xfEs/kvxJtFdHJe/PBIB8IExJ3mMgRtXK/QKNLqrd
0XnLT8/Sgkbk1Z30iyiQpMiiXnkNnTJNLPH9Rcn+1kL3SITcLQqpAufHekWAxHH9UgpBHMDD23XO
X7UaoBHCbCljAxw9+ghknEQmAu7YVqwTcPTwDUBNocPgYGnNv1k7UtMDWNwXMrdZ56fqdsTr5Mcr
tuelkvZnc8Ja+qmbSW3/NbMZxUJzKY8mMwj6ZpfLhzsjr7Z+xIOpXfFMCQ2ePAwKa0XbgZQ9y2yA
WAWLIfb0og+dn+A6jFHMlMcyki0c1YG324/YWFOdjq9jlPidxMMNefC9dkks2i7Lcwz9fwcVupHo
XeaAFpFVV7x+PEq8EXT5jUIaUWbqt9plkdCRJvjwloG7qa3ql/DL6wYeqorGli6EG0YZf2NUAHzs
iK5SinjOBy/FM/hk5soquxdlv4mIKPbkIyDiYls5iYwRMukBdVtmn1rejv5WVurk80SNUY5518jA
x/DfLF5DKMZdsX2zJz3yGpMA0Ep7zDiWlr/a+CDuH6F7ync6SEHMSyKzPI4yGPS4/Z3pKoMSDN6I
yhbp7FZWUrn62yCjFRsaNHQaHtVQmaFyDHAR2BDAbvOG1pHmdO0+eF5QUH5pWF5ORQQl7RWFJrdd
96721PGP+EwbLTfTX53z/LSD2Vgknj6dM2Zq2M5PQVTTsdd/p/DCv24uUx0PO6mTLM54NSTDAkR0
aOf35YMeX/+3VHoABZn6Oq/LGZYNoWTOm9SNqwgLjZfKUivnoImlTcLgo9PpFSGKNlH7cdoJdPBS
GRC5dgxxGHRCHtrNZvseLGCnXqxMgnt0HbQZzKmXltbv0nTzg8b0TgB/yxHOrBW9d/y+5snEj81G
/D44WqwaNG5cPFLcRzttMorcD2NgY3/Jt03xHY87WMAtIEJlzlFfebQn4vqKVmFSbJUqLL5Hmxoh
+a2N4mn/w1dDchBr3jPkCbBKIqH9vRjRYldOXpEssaVL9vzCmHsvQaqdVHdI+YFJqDH3y6w17VOU
I6msC2Y4MH/REs/YZlfCXrw+7MRFwa/KqRAU97u4Ym6icn9BxX9IJE/sMILElwkRnz3KCSM4yxXx
Bsw1NgIZaaeJJ2P9Npq4Q5weJKOAoBStEhkx8+/zpTF8t/xqC3TjGESCFCXT3vnDUZS28TIcVqFs
z6is9Z/HFlIa0/1nlXCOCpz+cLBFJzzhNgo0QaG2rCCJCrl8UHXz/n3wTOlWN7sk/QzRS1dDMqKX
UZeleiVMUBq66Sr9nu6L7Vp/X36z35vcFzIiJsuNg3PY7Nq5X2LklW52G6jbxkfniSOmmTgjQs3W
4Hbg3h2/S52FoCAGYkjqSl7e7jCfmQwQrGd1bXIb+NyjCnWZfhqTdtESC2NaUkksaEufvbftDV0W
qY4yTB15MlBnT+symOBm+YrEGGXrDYSCYkn1afvpO7MiDch04pgqeZO+d9RXWkzB6xGgiGCfleln
zcElcruiyLacqgXosjhJCyvGJ4EUBgs7MtuMdZnXg2V7tUnX9JnU9RlZcFz5fnHYqG+tMgHW6TZv
/JKuScKyz4Cq26nEaQHKZBfkAYCiaaXNa0D2qFR/f9ue0aDbEXdmVEXJjfTQzG7Jdy64dhWjvPBq
hDPyNB4SxVMwI6kqcpu2RjigYGBhz/AyWpPM9hZkz1yXkOMWBv9r2XdrpJHsDBaKhfIKMXG113Qr
1UBF8YcUCC6kSWFJ1eI0SECCtmXjs7MXmlZl0+5Z90QZlrZLSTLmjw44/EhTlC4NvAgfC1PLvpDQ
cspyu0nNVeJymkwhllFAtQobpTDjba2ehMjtnDqBdi8b5rRjy6zwT1hL9dY1v2OEVuu0jPo2gtOK
8Iv+Z1V3R68RnLzatz3JoxKjsreHx8bLO1n9GddRtvDBk8toI4J9TkAk2nti/2iyUMHUYAb0OSDF
J7lyqEvnkSa0OQ/cNWmoiB2Pktj2bauBYOjEBUkO16WnLBiN1c8rWk5peoe6+4hqHB39uRzfDh1B
1XWZH/mKSbIdNJVFpPmgIMP7loSw/VIys/Q9qSDOwu10HOAf0lez8NIkpcvOI+DmMW2RG7cazs/D
858q+Az6ooZH7VZXuQBE7SCC4m7eKmi9q83pF8vk5Ql9vGyjbPlnW5xfMMbofJYrvRCLHbDr6XP3
ji2tXbzNRLpOMGeilM7uy1t9g8niTpVSItC87csFwVSdaLRFczjvIXu2vQU+2gfx10fSFup3130J
JQ0xmqwhIKp+UgZqvrR20/rDwFjza4kOp1UcLN4OKgBOsQJA5nCtiVcMWijAzIACnfwwTSGXPW3X
XRJgO+8WNPpmbfn7AAWLPIxVZWbdXR0LzwO618Ytst0FOjkZdc983zpPsUcW7pE7ZRcz8wfK4WOT
SRcG3te4MFvpk6gA61ADwgzP7cMo4ptCDN/vHzb5eSxHMnoNAylS38ieIH0UEVwhW3ozTkdNVXEF
TdU2RXaUNegs3V4u/cu9zWTU59EsBmmIs2tGM/UGe8raBZufoLWv13Gykadr8IunUiSZaBXKSlu4
xMklLATXBwr7sQe2DeKWwkwcPuHnjk4v9B/QhOlDYz5ELALDwT+6W7gjY17Dfp5UNDYuZMI/OP6v
OLTC/ZCfwzxW/A7sL/iVS5gwr6TkXdFoXQjzyK5AKvHSnmZvt96sQWeFKDFd3CPC14sYm8lmy+L+
Pa3XSo9E76CRQPk9gmwuDruk9+/cc5nL+YwxbPuEPkPV/Aps+RCEFEVwrTRIr3NG0VoEWbiiZyPd
s5kupyXpveV01y6v05Uw+emeIyDBq4LRr2KXYuwl2eucU9nqWkE4+NaL4IC+DvnZCiQvpsYWoDy/
J9KpI5G4xGay5OTcWgGNWfLLRsq0rzoiLxvE9y7NZfQPHsYlW89qxwIkziSMJFpPZBs6PGjPmDbf
bUbml7xZ0708w5ERTsD8aE4mzfjX2HE2Rs5s0rJ9qsQE1ZyVR65xICs1l1DUhFfoAzGNXxk0wqpR
QfaQQQ1gsa1wywMmnCz50GTJlso0uHJEhvtJPSUfPZa5EfnUcdbrPyVBxJwDCsoop/p/5/kYf0dB
gcCk3pL2viGOrEW7rokx8FY4s1ayXEGTo86wbKjqYyOiyBDILVOvZgkffFmXF7zis61OQ7qs1Dec
y9eq+87M1Tzeq/jOLeUe3Kg3ioM6Tz+Gaa9dfTBHrmGRltAbUd1GmRGd4ILcVpO5MDLJhFSqfBOE
daUVM1+/Ukqu5y1uGpE/KvrmdEhEq8doiP6u2SPMt1QKp9Mn7xMq7issJ27UmWcN5YdJC1kHah0R
VOxJiJRNdDWBm5Lb3QdKt8b3HgcVnkiLQKh4zpZx/sABRUNyiqy4e5Qg85PE+X/gA3FVJwMDEzG3
n7UqIiugV2EINL/bnX6CC3UkU1rEVLUsmeU2/3HcVc/ePdfSm8e3PsTq60gVOf6UnZr9s/dEuvew
Pq6+95RPOQhJMtCYTnszasJmZ3L98M4BWmzkSjpGYsYn6GSW5zFc052M24e2Q44et7USNUNs+YpB
r/is6YLVo6RfrKMosshbwC2z7Xjp2e8Vym3Sf2MXyboGACBOPajDLEB9dzIYDwJwdp5CBgkX9ZsT
pmTgSKUbJByDtlh+LZr44DNS5q7vuzbS59cDGqHt0FOmL5tVirsevc0ZZh5Q1WvDeQ9n3aLMb0Xq
hd/eeutzt1zHSbxjaX66o2Ka35qC03ZWjo9QWDaUZ8pFScow+VyKGBPwyaeGW5LOUI6eN9ejD/gF
VfgS9QQUpDSBcYJQx5eA5PSSGzD5+q0w019ObhVsK6Lo3vzVKcbDm/X2+Sg9w3enTOJpnhFmeI71
UtmjDD2kz92f+uuMBFbgpKq3S9vyRn4mAbxNDNGJT+Qmgu2+qHv1Mw3KmZr7VfJrE8ZzgOM8BosT
VX69Ypo0KG5mabPD1SYjlrdUVBtZfZjcsUAwjzcWYRRjdf4zac2SOiWbgcuVWwTuw/0Zk/5Nb78X
LjLYAZT12coStT8Cr1ewccsSwONj7VSm/fWEa+K/1rRzGUWH+uCnsl2D0dGB2+vE7/NZV/MmykjO
AgZwwCSbbZTnbnVEnCXIlNiPnDQLs/vX2dBW6jnWUeXdsX+okhKYNwUow5bftJ2sSrjYhEO0uv0d
B6m/yj2kqKwFQv187Ofq9Q/YzP7ZskgS5kFQq1ezS8JMH9R3IxxUgOHKdUS8NcbZbp8kV7ed6z6t
XmFl56q4UZFnpic8NY904+fJkPOFCqPuSsLIuv/4gztVGjauQtQGFHW9XGAHw2bvP773BSQMdYAn
l/74N4bIufrlkLS3cgz3kYbMs2kr9roIcHadOjnTOUKc6Dh7kCTo4FyQQ8xcEi2bA3q/wm0ulnZc
dCv0qgh6Fnt/yA3UKYtHgqAwOpql/vM9T2YbxeBkuPgUE694GzL0N4c0XNdmYGN2cuVlx5kLqt8I
n/wd3CB7Degv3Ivn68ptqBucV8DG1yamJTSeSNCJztzmLuYswTRBTogm60S1TxuWr0z4dDiyvl2N
H8/7q48iVPY/OrydCMtC7i5VlHZ0zyAQfCfLmy2H9JQb8B4M4SYFEXHMyvXdjEynQIJZn1gd6Rcf
V2XC+Lw2pt+dCi6JhdKssXx7fl7lFr0bqNQ3fU+6jEOjE3kUoh5QpEhztp+ot8ejLu7k1zkSYrmQ
wNk/QcCoK4ZUpiWdkUttoei4wG0q2A3QpYM0TnrnEgFmoyBRn96GT2MyvPWcz2n5BQvp1VzPLu+b
sOVht2rqtVtAbPdciI/DA5LYrqnZc3Rc3a1BskFT0DR6O8GkaFqZtPhp8d/EbJ994XmrCQh7K2iD
ZqsIBK6eYnR5m3YrP5xUyV/dlrwjnm9D0F/gwHS9OVT1YVCIfzgR16sn5FMNI5nFX0vvWiCDEqR8
VJeRSo20tAX3EAz/JBGi2EcdqBcxY3KZj8hP8nZjtfCL6wtFy5lumZ3Zq98ShejH7S0/gnLTryap
XqWHKYJLx46BkNxDmlBXSRj4BLEbvjWK/L3jH4pENavU8UVL6JOqp4ujjsFFxjEW8B9PI/+tuTDf
kVGmbMaFC84W9QT8H3Cq3fEai1wSoWL5xXH0icWyaVsGpjJpgihFXrztHEaqj5FtaExpAIutHWWS
UvLoDZN+mqyO+nCcKiAXqj8bOD9xAZaFKFTV3QdDf2jzq15ES0macvpV0Xj8YLdCS6JSUUJWM4sE
u8s+2P1yWpk1ZuSbb05yvDa47caANHh6vJP/yg56QK0aVQdtNsFTcGe6N/ohfSd1HxI3ovK4BaLp
nA7j6J74rtwywZyrLHlzE6/ETPS8A9pNZPHIWQHnGbcK/KwyweQQSQlKGnhNODsaEaGOixiZ2Xp+
GsaKtT1WjImVjK69IwZ6LL3ZV05DhYEDBrCzwvn4byP+xH0veudOnbnCDF2L4HZ/V+NOjgNVJqw7
nMs25T4pE2twmrF9Qa7uo6B5szP0WjP1ADSwO3+V2CQN8XvKXk+wKW60UddK60fXhVhhYq+qzTx8
63j4lQ3IG+wabYBG5q/dxvHibiH+w66eTp1eh66lBbRQ5V4nyrvSI+i0cLGNHmOr95cfUmH6dpYJ
091A07Jgu5Sa//TCGcGP9Q8BRD8Y8LAOCYp5XmqlkVr+oQlULHWhlh4nxEtKfi7Abi8cgB6frc2Y
lTjfqBfkZj3rCjFw4tSTuKrbeqVYBN94BrEEbd2y76PpoPfIPUfbv28BO4FWRhC24RSE/qGqqD4x
uTyOi3z7vzx1zfdWqI+9A8Ph0FQIi9U+x/wPZ6/fZs0eB1eVixI/69NnGXPHc3T5VcaSxJSn2DyU
8OtZu7QE/DGmmfIMyygEt3wGCfRTeqVbw984dli/SYCAsYjlj15e/QNbU1dnBKqPzcDafYlQqLp1
ouSALk6HEZ5lNrEKdyECYK9lN6/dbdjaXbfrUniZ9dDoiaMghgU+k1cHZq3TaMvwksuz0/qSIwg3
U+xV3C3vtVyhfKxRtr9NvwFjf7yPF4K1lg9i5p2XzQcbNOhAWzV6aKqWTjsCo14d3wEwVRgRRa8M
THKoypIvGX4P+YYVnSOfqvM2iM+gFrwT9bcJzfeCkGeBKxajVAVH+Q/+mYKtAq6nfI8WmwY+NVuo
j9/gWHwN8fwFU8jS+FBbbdeGNiSN91zqST0D+OuQ8wavZKDOn1gjKUMwiUJ9FxTdZiIo1BTrpxna
46c7PMyvlQy0xT53iJxRy3P7BLyz04eD15JVNycMC+elgKFFyf4U/7eyboK/VMkILLyY5u6jdUNy
w7fOSqKA14ad/ETF9ZeE3hAYLHYWNPf7Q5H3HJnILLSlLWGdumAaqg+40jJVtypZi7qMA7DlJEI4
5X+RBNFNBZImqrhjIGBp2Dsj6AiuWvdv15Hj7Gl7UxYQwL4i8O8lWQMz0zOhWLZWd9YwXtuNm384
tSXTAe7e/WkoIIr5wtYyrfES8FXa2kFI7so6TuhVcZoQ41347yZH5v0ArCMMsek+pZ1VdMWdfwV0
FDyUrPuRLKvgcZQSI3JQ+rNmtaEOav3SnvWUllhtupKOI7gMa+OJ8sjMNgBahxScU1/eLsHbrg8x
11KHVFSsiMJaxgf1hG/rEtIaeBghYzOMTvvkkMM6AXdQU3mvNrxEt94CjYpqEUmpg5S1qFxjwrTK
BqWHieA7ZN32wObtuoSQ04YrYBYEoU1OuHBs+t3xhkr3Ezj2QHBGMMY84GW9MTw3Yf6ced6QMFHJ
tiwjUK2XaTbWbvt00WyB+21uREvMnngXOHXY6C0a0+y2dNmJ1/raCQQZj78ZHdMuccNP0LPK7+Jk
NglCNYHNbYHJlL78JmDGErCvFX6ImvqoF7hKSxNWJ2JsyIMj8VdDO9mgWuREbRSzg0AdBqZ0uFXf
oDMmU57KZ0WQJRv2joat0ODV26fQpbWuL7LE2Ww1P6oOt7Uf1gCvz9bn/fL6JbQxpGQXoLPU/pCB
CbqlKScG7F9KZhqPnO9PJbi2gdW1vku7dXypsEcJvRcQw/RsxrfoDBS9voel019IeCgmJHKzyz1m
AvMMWvi/Oj2HMVu3wGNuPAFwMVCMsuXmMWbGCiAn/2j/jhLlQIpSUreTGk0ESDin3RGnOulkKzYU
83M6oQD87nIBDVuqEng3zOtAq8oQQWMugpJii5VKV9HJL078so3rvHN5gkZPcA7lfrcTGkv/l82M
s+oWzRJxwKemwhu6o3t/8KWfSrt2cqoK+7FGW+QrIK8BF+QR7IlYqCQftgcIOj1MkVsjELhZU/Bt
45sNSdcl/grmYxTKc99HZRfa5FoQrTD4WrI9NIJhLdcWSHlAisBgucRl1M0MqTzWEaSkKzD/d+3B
mzo1Ppw5NWccm+FxNYAWmrk/dKM00mCPfjeYogIAughmoJToF/+W8YuZEAzTZozwo7NXqkiH8bMp
/9ITdUiVEfsj0jM8gWwTTWIqPRNkgzbO34E2PIu9oHuGW0o1WStts/ES/1+LI47LEjeIChATLWjb
jullfxVGEPM2HxkC/+l9NNPzoURwz3AsC7jav/aajMpr8MaSVtnWJzcPTsr/U4VkMMFrZBAVKrNA
KAyXy5yoUQCmq3uLj8qtwIadaZv1OjOxGZfUUprXKVgXt7vFtTVWDC6UGtn0yTnXirIIwqwuFrOr
xqiIoEXX+LOi3DwGdRvWFBr7mavqTNGciuVVS+KHhC1Dw4CJzXOeJvie62AHgoRbLyvpGeeOZ1c7
n768n1l+IW0yMcKnix0eXZd2g7RbIL01pxseZ8DZQUcAF1XXkj0nWNoHF5WJ7JzW14839pcOB9x2
vnov221w/Dx0YC5IWVIFS6ppoQYrXUMg+wHLHTbJYpe8ksJKAdreTEWGvIwtH4aizJfnW2FY+9WL
Pw524sWynArwL4S8Iv9sWvpev/FM+UX31QXnachhs0szuOB4TKKKbCGtuKpzFWHexMR+P7Am/urj
2WnMCHNGQf7o8Db7oeqrno8sxF3E1aC0xszxRibNHATarA9ak2NReq1DU0YFswhZ8vLTW9cMujuF
MCGbVAC9EKJ3mX+WZucpDWHwrXA/4tp9bt+mkQsWMcJKSYqXzV3r2PALONHDyc+MfcgRw+6GgOqj
yz6QZoJrXC2Zw5F4BxgPfZnosc29KcxkdrGpcuYaWjCQvVBsGRxQ9+FHzLd3/pf7J1qICw7w27JW
pi6o3TJ+ns5W1R2dY/tWLGD/+jOjnb+UC6nTxDVx6hXLR3f+chffLt6HWbm/VuH2z+UOUxelfmd1
5pVzY0/VBiDwuICCA8YYMofNMQn5C4+0jRjmK61qYiVY7fCJVv8zClQsZYBmGbQDKaMKg6JSC7/c
BuS+JDJfD/g5XbFs1fKkDIgW19wqFHKZf0+YSNCq3rkkgCzDNWSg7TJanlHet+DcSeXiEM4uWS3X
Gvoxy4z0SLdw/554e0sHKa0xifDZuBPrRh0tJ+EDMT36vK2BK7fH/BvzUc5v+S85EGQVgJnphWO1
1alTGOjCeQ5LBD8tjr/yEpoHBPw5ZGcjr8YyECChI3tH6nwaRZAOrnGgOFM9cJ6NAcR7fcgK6xI9
Hz61BAuuCv3RD7z47Q1BwtGU2PX3XWmdBxG0whmX0T2Dl9nQY7m53LpfnikoTlBMrsfWbWgH84jA
7O0YfvZXSMmiGvRc7kpN/vUttsdfrjppKCiB1P39vpkz70GgbKShChQtfgUhSMuviQMVJS4iTvD9
QnuhDn88j0TSltps9FN20vnfGviFzrh8Bj1Wp2lw222PXhSigEWa9Zp0jKXTlggjNyj1r64miZoE
MFA0tsqNFQeDHPA6BeuNksibWPlNH3lQuJ/1ndTlnlAldPhQOTjcnMLcZZSvqal5m2waOIuWqAaU
RGOsbBJ8e1borcV/pEfV02a2x83hX6aQ0+ZjQV/MS/jnCF7wrGXg5ux8uNVgQyf/rgpsliIbnjiF
Siolwf76IFSk8WcdC2+Z2uQinqyyaWGGbyshjmtYdpaQQla+lsMKhkv3nfCqxNlhFMVjqcPLA7ea
Pln2cqBOFKF81mSsqYW7XPD9pXU65wuZJSPwo6p/hD5BEKPjdY2t2z+qs5viD/77zwBRcRNWWt8+
QW4bQsNgm4gFVN/o2sMxSomldKTQ4QRsLuWTi1fJRTNh1SLnn1LIUZpdzNw8jfMO33Hjt6zKfBa+
pf/xGCWiSllqiud0kfyHE2fxOsF2pRlfhPj3cwd8N6U/FPOQTAO48kUfzoaxbcfXbaFlhQA9P1A2
u2B3dvncLGHcN9p0nDC/xeVnnFs22N1O+KUJmsabFbzHC+sBP/g7U3G9/bSl2lH071A92RZubxS9
5TI+QNw9AihUxq1H7l0eEmIeFQAbAStDf8ujiB1Rl8WMS5rUD6WlpCBwJsePPx1f4KcqadFUrvwR
8/yAqREl3IlODt0X+mWPJGKgCdQKfPCuIwAj+zwwjx+MkKe2NSYgeZ4L7M5rjGUixvgci6WOyx8l
mvYjBBr+fwthMIxwM3NySdG1JFVd1fz/8dchW1qpAaf3tBId6Rof7ZRWRm33T+eW/UdMRTtYpQXl
nlU7Pd4Z4Q6Gb4djM/tn4e0Mnnb5TG/v5+feBAkP0zO/f4GSFN/AuHMS3x/xJFd4Yp8So3gMPvGi
8LUUNDUDgfpjJDBoF0JFcyWiqoOWB5HmCcyYUSq1gGZaHw3Ou5pq0Ci2PYb+hNLl+7uHMejH94vd
094TBib5RqwVmeUhxVB359XkasDFJvqp2pOVZ/+d6YdkV1BkFFp3TRpSAXRje0CLOFqKAbYSbFBy
+BFT5XpthU+OZ+1ufFb3YjgJiNo18DjTttPoGODJlYNIM91nen16iYSvA2ufPiV1gC/QC91ObEwI
0yRDNpXx1Xi1KD1/pVeOeLG2A7eKT9J0xMCRtQimkYf9SY1mQ+e67DUunyLylbLdsVzxpijtqgDP
cOSY48Gn85nrwy7kBaX+HGQNNzpGTC3HJHPqahVkMCEPRwuBaj/sH2+lGnwesg+83D0Tc4GgKmra
P765WvBVFI7+safvFtgFAs0YJmIj6Bq/3iKrNcLzj6P/VyQJlJm6D2z/SIUiG6CJrmSfKDmFWZXl
qGxk/N5Vya0iAIeoFp7GZOFmXESJNY85CbpaK5nkqrIj61CYsZN35P0wWAlxnGAbTg4I1cEPSQdg
hllCx7osH3JJYGen0Yb4NzePw9btT51mHquzq5WMdHnOiOavII3MHQnaG9J0oix+EDrPRe1DZaoD
S6MaZiUt2xdin7zawmw6iCLsz64jckfB8tS/a/EiE6l4WfISQPJX3EMLpcAAQTAkN7l3iHdyPaj5
Ww4MCXrZb2R6/KeFw8qrsZk6/qByov2MOsvkORylZ3+YUQ0+DEEv/TJZihwOZFb83fqIS5RvurZQ
bn3wO5AQv5TOcnzRyLRzjh3ersuLWBZTMEKcJIILDZtN65vXV1GNX9KdpgVskN7GhkwHUVIhNiz5
Y7ZBiSc8T9Oh73JL4/XZhgUyeiQ9Mz1pyTxLKgRsB8iXK/vJHoI3nJCELWq1e10P1FSisQksqLSS
h+zuxgZmTw6uFOUQ9M9IIzP9KATb8+x61wSGYtp29XrdK8HnPHklHevNHiS/rljYehEpHKoXr2Kt
NZg8jvSW7ROwOd9W9BCfqG3MFk9z0mEuWN/xVZNtRCB3w4m0UuFBBo8pALkOttOThDbxVGp/8bQR
Gpr3pwqM8K1wStxm+LJxD1Fpx5UmsorxYaPUjmJazpUnPTVQPwOuCFSl5A1wBDUoIfMeU3DpfiOf
pkz93R/XsdCjq8aROxMLowQhWF/4cqWSCOSQWPoxyNhvOYeB+wteSBa40tCGbJ0BtCNbLwJQ7g7x
x3tA0tnlqFNKUpITbQ5OqrOorXrilXJa+AqCYECEXCqSFa2idDYDzAPMabDP+M83rPUiJaJSsbdt
zhAJLwzAlYyVMh/jfUBDnGOlmklHwrPYX83j85g6pAPfrJnLAVXS+e9TneRK08XgPm1wVf5VhQUU
XqqzzvVDwmGIi0Ywec0ifoiQLupw/dSAe9hI8MBPoNYAz+z2r/oXMCnWFJeoRzQ8AhZQfwLydCb9
tRwYjOEOJ6MYSWvum6d+wALtnQfFHR7VE7MwIobmPRf83r9N+sWTG/sj1rdhi4bVXPq3xeM2XbOf
aEclPZ4XyFThGk2BrTdl18kxJrFsXWwLz0THPHYPRIwjuhLiAxclbNFmE0e1ydfMNxLwLI0hQxdy
yPLnmjzhmYKGLv0+U9LodzteRTUFXllHD59oSbfEPcpi5YcGoTeJ2PebS/srkhUH2zX9zF1TIeKX
a7gcYm7keJ71Ytm4THlRhjLhGppXoMeR8cfbU/iHfCiUhAOG6Z3o3xmXm4W7tb//CHAr9YsMI1QF
kc9lzM5VnrRCZXEMIJBzZBQheeXY74bgR2mKJIeVU/CWTsn2PM6kFTwlrwWzUVcPn2dBWGCSp26j
r2O2CQRaVEYjdISjyxJxHXRYCWn0tKvEY3FsHMSAjIx87SgUaplBNLyIVdcoUj1YFQJ+ItZZLWBq
rYlMpm3JSrMrp8uRgxmCcirYWEq9BlFeXmzYatePEOuoJ0gAUlI9UV4q+dxoMvE0WrtYxvCiwo8j
vV0lnjpvCc/Y4iJwUY/XTuqLVLM995hbhWYO5xmQfKeeoZq8wKHJSUC4nB35XimL5mtfBmcoACZi
BY0PlwJCmT1fCYdGmgDVNvWRR5Zni37KsHsm3lTFREUfHPU/qbXjM6wy39UPEKxoe6eWwrW/X8pi
qRXly5Nh7jAjWeaVAOK2r07VEVARke/XemUp6zecGlSBnKMbvnrg4iNgN5D69Q8cn/lhbjqqKlvt
gyxNkRLCuFvdlb4UGXzb6F9cFlbJi/FPrI0nQHlHKV/b8g83uH1n9Zs0eRdWNSidAcZF9Tlqnp6X
Mxi1MxWvreQiTeB+f4QGxcW1iora5blZnFliLTYU8qnrX/gf4DvpLilZj84fI7NNkaGAP0JRfCZ2
M96ERFEaBVSCnPBws8S0XUAtP/1hBhAsDEKCApDrgs4mdT1J2EfW10dvunk/ntUyX3kLK7ZWAlHl
vyQzWjHSXId3dGmMm8JkDmv9oi5fI1M/byrUnctEmgDBWQK4nTR4M21FpCF2b/f+0F+yRRK30Ic3
kAv29V0Z1Y8ziaLxO/UsYyyW09opp+WYxRtVC1vQRaQKVH3dBKzh94Fgd3hwwzKWladHJtuuGDVQ
//CU/MM6vg0N8weLShGavKqCPev++PrtrxwEiaWKUAUUbqqmlSm2HxyyBqCMkTas1vPQvYEm8EMW
HLzNxP0a/upLsEU6zWFUW20OIXPff4P5ZLv2jDhLLO/4+VMgjcdIz3bmFdRLg7iRU60mXoBF9gMj
+bqlAMiDUsnAT6X0QychEuDay2FKnvJDPyFMT9L2f4itvTcYBcquRqjd+r/GyyIn/9M3tdzTMjBZ
QeVoMD4Vch3Y1kAYbh7s4mxliPPIrzzyqAdamMOPscLSsTYUg3/ITOhbsn217eU9KzQWjJP19ka7
dGVEISzOoFQiWyRitZNV3vdzv9T8YmrJ0tVpvMLtfnbB5R66UMD5cC8GKAx7NdGxkkyNCWeqdcwf
FRLVOkx+VVfgMKzWy7A6Zw2aZ/0vqwQgHdLmshzrWjbHNfr+ERWhhbVxafgaLYzC+fXlxBe6CwUN
IKEMRMadqp4N5EtG+SfrimqLztLL+3w8rK7xi/MlYEcwLc9wSiMsv9JDpob/hY/pkpBXKGWxqRN/
Awq08iVg3NQ5Vtr72wXkGRBRAni6IwGP/ivLgMvjYhsAHkTfetTo+bGW/P+rNA9alMkRlrXjoS7v
ERqnaTOBKy5Y1daiHIflFTOhhfu+3xORGSs4iXpiRxoU0fZL4EFMvPLTL0v3yU982+ogKAs3tRZ5
JurgpREMW5AFHkImabDTPZmi1lclpFUp8A3aybnqwaArmcF5CyoLjhIs64CMlJ5ALNAjPAzLm9Aq
DKzWVjvcvdHzZyjWUR94VO+4iG/wzkJfv8nYJt55gybzOZ3k9rWZT/fk5ZmqKWbgRVDuGNTFbboO
/PFgmRfxIqkAncFlYM8yHSICLxob5a5vsOBkxcaiiP1PvFoG6RLT3Fd3yBJYZJr96fVLorO3qNiO
TfFthsqb1HalH8EDrDPHdSN3MK9N7uoFEYA8iIGEWAWgej6h0alP26RZ3CH6OecA7qnlzomQ1quM
lcjEzj6oQDZTfGywntQ/fJySn/JNcZMnlQSubMG0AeHwtRcK/WPxyq5KciB9UkiN/An111/17fys
cfl9TVbmQMHiRff/x/Y4CTmX0ihUnq1vuBypHOo8Ozvc54xQzO8fMwyYCOiytyUAjYXJ1s48Or3e
9b8wCFjoeH3Ddy61nfA+Lp5UXupIzpincT31txa3EL56ZUPiE52OVql6dRDuJZ/22MsfsEsNBkxV
LHDFmEO20ZRI2a/d9TGZi+tzbEzD5WbFXpN3eBxULBoecO5USVZRCtUQHmUDSeVplpDbn/7LZ0F6
37eaqMDulzlMk5e2nsD9A4DI85rT3PzDdRseAiu7lWbCtqsvzYo0h+3rTh21MUAXS5Lfopj+EBgx
DTc3OEzOz/7GaSB+nS5eGlaE++ZGV3gjdTOjBwwaA798xF6ngD5WDKmk6ozdCQt9IzvM0aSZel/9
WxDxQmL3+3HBiTMYaQFsPYRutbqP99X0QgzV09a3GNx6HKAvqBkKtx4i6+RNd457Fi5oSFCO1a9j
iFmYy5PFX1qPp9v/geI33iLKJCE+g2eRL/6X2oLKB5zwumobGa1RwAgyIsq//+0/EA4NFN5zlmOx
uRxx6W0RUxy3Gehg9B20l7OBIgvCZuZOnSNHlqDU11iYlSCC2Ctl8JU9ehc3d+hBjInaMAcy6Zoi
Mf1flN4696zejMr2Z8Rm6uNiGaQ6SH3tjYONqP3ziMr2vm9Boq3zgf2Qy19fNu74e5sa0r2GBDy+
KdnzgS3fH6RiLOvbTr8ul8DMcTig3PwvzLXj/Xj013lz85vCqRTnZt6KfcVr0Lws4qXieDc0m+0k
hlUvmKk6n1I4dKeyYx4u/ITdLvB01B4ek8kh3CwvfMYb+3TtG8n/H7xoNrfcTbhJPKYBmT1wt1qo
AGgxMb/UkkY75/SywYhLVaktfL24V7o04C8o4pN65WF/dY4cL+XnSdZ6wVp8vlOcDVeI3BcwRcWj
Aei5cvkxWutOD1aUgkmdNYbtqdEHNKlhdBnNpIGSRQWANZpmHw7lrV0Hy/qauPuLfAjQaetcd6MD
peOmv88SkacMeAy/rAUV565BU0Z49WjD9uRNRktB2OyVnEjCCnQge13d2mPuVGlqIte8ew34jMAR
JzZXl5MSqmU9va5Qosrr6xB7Amm/KzSWbVOYQk8by4JeXPALUhB9EHsuUjMsVkWN51EWhHcnwOKs
j8uqITcgIytDaHPUB1nKvWHN1cmtUHqnWrzWryo2X7LCcIgEmqrbpVb+XceWfXFErW+9zEKoZsY3
Z381y61eNYFaJuu294++y4uxiWRQAC9RyBKVKAJPZeBOFRDtNSapm6z3hJxZEP5nxpI0l8gNQjTB
Y2uy9PYpktuRTRegln38rKvwPgMy77oFCOWiXpNoQDs3jCnghf2PabKwh/YQA2IlbVZNgOWeON4I
CsJdG5+lO3MOnSGi+O+j4qSJJmNij/XObZW6E7/yFO0bDZEB5xzPlgK7v2RZTEIBmTS72bHw7xKu
qcEhKlZInzzkZWuqTkG6fZgnnp7xDCX7onQKPSDTaVuaAV58lMST3MLRKARJUIgghU3mJYW5XLwh
xJ+1VF8cUbFoTglT03fI2goC9KR3db8sw64XHZxgkF44hg0xaQAgVxeH6TVBoYcejZXAcGYGuPc3
NvVH1ly+48BL12eJXOZMcXl2PCqOf0ljp0/1nWbsfUqkKi8Cbr9dEjOxukPjlPfUTJd8i5oIUY5H
zZG0/il1O5yHl6CmApdFzab9VBbZ3abTKIWymEbXlsSq9jQj1OPFER/WkGadgY9b2FF3OeWC5YlZ
ElsZsw0Mufa3OTODagKYLS3LM3+wSGRZV0ucQK/ZY3yd44LPAxJg3j2kIQfflsFuKoqr3cxTBFBB
b4/qJo9nMQVeEC2qE3xByN/1Wg/wD1VrqArXEkty9eKN2DDoEz3bBN6aMKHZTHuR2NYSJqMQaB7K
RhotuLBZ0dgOVQqaSs5wLOkt0bNR2/1LFHdVqLh84xmYfCbE7zEwaLEmFBqcjajk/1wbsVgwzLyv
1hhl6VbXj9X7h0dJjDnbmsz2QdWRRqK+4HgNEKBPuEKInRUGgHFVckRjiCeG5mvMzwE/ad34edjn
JjPkcb3wBMD4IK89hyParsbyR/InX7HzJA7roUI5tPWvP8jZyhTFrvUak4uxe89UXMt19viEXITA
g6P+9bg6I9CaJeeRophs+6tEBHNRJHK9rDQgaLxV9oAX9YHmcVmuVgiGqsoqGCS0ds5Bqn8OsDmw
16UOqbKPyBBBUI7WrAHrtBaIUMp6zfk9h29HaP5dnHVR65YNYELh0XvYtCro8ZzsXTUuROZ/36To
41YsVQaT46D7c7fj5du3bNFuo+xjFxPpqwK08KsYbmrscRDJO7Llp4SYME+IVycw1/AbmTZpQa39
oKBBF93CyFxNcx2kucIvciVj92r9jfUstIJ2kgQmvX9wNlbJ6vcyhpItShlDO3sfhuijck/gqkRh
YTittDdxkGGgAVerAxIvI+bYf6i7u5Ho+/Ca+nnfKt0hcjGMsaOmFBUJsKt0q8QOTWVgtKdmLQnK
pluu6EbijN1hR/ATy0jpNp9PGTheZV5j/mzR5pxI1wz45fGVtI1y1Qjl75fr3ibyWI//qtnJNy2Y
23UXkj/hcDcU/aw8ay95ThuLksAYl0YtmeQkh9/LbAfvtaTsJtZBj4vofTy+t6kkEAalm1pVHwf5
bUQNRUeIsSgOuRiT3pRf/rYXMwDKZEm8slwwoTrxZqISQbQ04EXVEv1ivly66qgLctJ3srWY8LEe
fB0IiyluoWRWWxxw28xcZkeAkStHMb/A+84qRgDt/ZIhOI3CMDKJV7OtiZjgNgy0eYvEjfRE077/
HlSOcMVaH1YwFQy4qFDG6Zz1I9jm9WODgQOpmKTAw3AmyCUJOKzILQUfzIhPfkdAI9UPGtzJO8/I
2Di0VdUOICWduxBtwkoSVtLO6NQGgv4hYw6kaXkA+ZBb8l7/HhFHsnJWjyuEcyKf2hBF4Kt6g/ok
bE9luew4dCfBZn4GkHjy1ru3pxwALglVDdsmoYOja+CG8QLuP7pQ0gEhfrwknLSrMK0c/MSFliDC
gwMa+KpFlYrkqFbSjEhYkXsTsQkK/I8C2c5dakSjpNQtf1u7UTwHe1hmP4Hi8wHrjkJtR8zA0Fh5
TiykC/G/CRE520nb03MQ7sO92yegigiI8gT0/NBCY/53O8J5EN/UvkQeAY4YuDODtwHYmQt6lAZn
8TaP4bXtVMCcggoPlfbAGHZDson9ozl6dUBmOhkYjqA6Qa/fkS4K02RZpFF136a3ZsAJ+90EASxw
oxny4HEjwaDUoHse8vSUUoLZyM0FJ+8r2SRqUC4Ksv6n/qxK5jh3GxJbPe60kjwHkcxsSKoK2JHt
KaodUgVhjZydbKPfhX3RQLoaNeSJkMwVd5+2Ju1j0CM9Fg46WpbOcuDHWLK858XLqoeIrZrTA90X
mwhE50L+jaljesEkwqJnyhQCITtHeQ4XnO1axW12vm9h1Boc931zwLHae33pOEFwmmZTrZJRuBWx
CKWMubfbp/6pgBNLNu5ZMroxC2zLP1fku1WXutiUCRWNc4adq9SY0RI/vOsFoWXpUG4xHPlKoJA5
Glw5foFHQCzqPkp6IqvukMr6s3PT55IUcdTefR68TKWKV8bfh3LfXDiVmmfolUIeKYAxxWCVI5NF
aoYTQhHtVumPnc23N20I/4xYoz6s9SYuRiMQeCYm9FlkJhrCRhQvyEe/yq5ihDMyyBX4vuyfpSIq
VZN/iV2mAh0q7Vv5l/TnXn1kr9PSW3m/zajuNFXF2cuUUcNUbDTCiqSXS1/0+UkgTdp015tvJ0fz
i8T9OIDunkIxG1T5UhTccsyQsztK+UNiaTHzD1Zp3vnRzaKv3tbpKwtgZLCpwxNutVgUrKFt+zqV
m6ivJb+s5Hf/q0WcbYQmOu0Zzysd4SSHaXEr1RhBoZfLbv2pIoti/DHiycOzFOsHn1tc15gkWeiZ
0jZtHb/DsGYwy7+mytBMzY6kHJfS1+o9WRZecPpqooQf5RhKFI/THdfc22JnrT/QhuGrYUWMSY/v
BO64T39lpmjkgJeyZGHH5mrYvV43QcYSvUK4/gIHYgmKE9iTnvQCLG1/M2OUTP46sQg4lxkCvNl6
b8aez+QSeoLnbMXYvzlWcnZ2+BClBWbWrJf5NZ4kUhr0wO9WXvT4aQzIDrre7W8M059k2i1BAD0h
MwAoN71BK+BLqec/yXZv7XPOgaqoaPixD2G7Bhm1f+KfUj9Mwr2h8EAbHh9kME9NhEIaNR7dSpCF
Ut21A1B4WwCQPwVNCioZOBRqPd4KHPTjswgMqKoFGCcYQMA5Bnis+NlcTb1PIrq62Vhnp24KUDWN
VrZAjj1cHMR5ukS/eEGfkAB7/zY/o9soBBanS0KDKzcIWEhuHp+wnGEnGK5qXNgsyxzca7T0mn6/
9kIXg9f8uRasfPN3OD34kGG1qZuCcmI5/L79EPiqJClOeWAigZAwc6CX6gONTaBzIU/RN2V1SLxD
Kxa4jsMFKgrIV5v94b94J2VxdAbH0oDdSCjANz+8xUoh+TGOIl8UlGYJ2f7euAU1D5qV4uByfTyq
bLCbzbn3wlU1FWcg377NgqWX1V3v3xfabvKYvsfeTlafxcbQRUquPVsMjE11u5mha4acSgt3qj2g
MATz6DQEqMhrZqK/zVUtq7S2/hGb5mGEhmC+QXBgbY2jpfK31T4S1lHJcJ1tEJTUJYJpN1Lxw/un
KLg7te+ti85BmDoumsSlzTqIfUM1aC9IHPZ4iYo36tIKLEhzkaGAwqbO7+/JLZSg5OclDEF7Pqcb
Wk+glHkiP2WyrRs6exF0fSkzDuN+EYJ8iQtRlKUzT7+5eL9VMK4wEA1n9TeccRhlPF2adtMhOGa7
DeMk+UwAT4gSgQZxefaKl1NU+0HZYp3AhctqeqF27eAYaNXFp4V5j2sFr8NhEtK96UO56GPeAIba
fNPgVjiOsTaMu78mVjFFrdYjCdz0uIDhcUMMfBpQ7MDF1EPIdm4c4Dd7rqCpmTjMkXNd9Zza3I1V
bDgq8mSRBNxDG98phg4RUce5RVqiO1Bo9qHJcaMQLtf3jG86y/13jIP5RVc3uN6ko8n056LFN6E2
scCGSixioUhoX3HBAuIWClj2Kv35nfiB9VSTgJT6KjkXg/WVN6hG2YVYHXyTBCGkg6L8TuDFO2TE
A2FMl6WigFnb0LiKNpJ6MqDzb/mOrsGcETMtagtz/WcbUlb4lhRbdfPk0IE0gsg9Y+qcuyGINI/X
JcUyvZu1/rYE9FQFjYEp22r5BRDLgYrpdMaDz0sYG5+bT313jhCmyDKlgjdPNw56MUpQ03NhZCOg
BFaAwGobz993hGrKQy26ZzjtxJ10J5ysTZyILMrTHlsofdD1uAB3/MBsm9sY4FMpWN3/dUEJlcA8
uQ16kAOf726J75+ZitBB9StV3BPyfIt1o2b5/5hCz9lpMn3MdQhVdC8dsdpKm/sER2dVRv812Ris
yT1XO7UJm3VuRcxd9u2nmR0zR8prUsLnHlb0eNtedYgMNtil1KDskjmn2Gc6wAz6/B6TMFd47LJZ
F0dQkK6ItJSsh72IbhmG7FoLcjXHKiXqhnZKO1UIrMKrnHHJewahCHIFAtd/zcSGCdT5TU4MMCX2
hs32qsm+0U3+zKMTg/QEJ87hxxzu3ShiZqzKrZTqg3N4KIb+BFKNMm/Wyd6cSlU9IsKn8jsuAKbc
+NT0bw2t5loYyJ0TQ4YEAVyqzDCBLqS8TJkX1Bk2nOpamf9ZVh7gMzB+8kdzEOIY//gKTmMt17yu
Aaomns0GOXIYCLszsRcgyMgUHY2IwQQl23E9CqRGK8Z1TSTckg4t1GWrwaHiXB9FSlj3UenzLimR
GZUI0/dFepjDLERTgwug/cMa4MnoCvx0gBOTPkdqTSh7oUHoyq2vKplTBnNgeVdDOqoj6r3WOVHh
eMmuYYHnYsQgXZ1RMLjs74moTXg4Y0vd6CVSj208R00z3OeDcdVscA7bEjZPIcJxzRoFGFz6k9R4
Mu18ieuvxdoVTu8KCjTRN7f3c7mUmOt95B+/EVyn98C90eRtuE3Cd4R4vexUiYbHINhHGylTJDRP
WvOM1t5hOyqP2mM9Wz4AxcCafP4v3IusWzVBCrH2qtD1gEaz7kEukapBy80TmoH6dJSBkNPhLWSi
QASb8D6CPtkv0DoT6EId2ajzY8oc3ZVbgVqxMSmS3PIR0X2xgLnRPq8Q4RNw+0a00emAZaF9mFbZ
FR9QIllnhdoFu3PluJMjGaeANDOO5PpLaWa9u130//FU6f79HBS9M7Kw7n5TsBBdUOl6wK6cVlUW
WFUuhi9E7C7NZiEeI54UNCLu0J+pfI8f51IvW7fTWyMOPHwviixZM5RRCkGCRhcMFxDzJ9+WM3Qs
2RUuKwgKeFUO0obv4GIyxGaAmfRMoMRJ5I8LcL+S8BMU57d9tCt1AgdrHg2GXhPyuvJAZcsVVB/N
oYn4x+bs6MSat+FAb6fbFSiO8kHLuNexwAvecO6pkT7KQ1wqGyUvKuQtIBdq+tO2mkg1dzFfkVQB
0twY8Ge6QNUYrY/ywOmoK4M2smGRQW1oxgQTHv+skVRUg50plgGmzdBgwJWvk+mF7tma0xcuuGCl
5EQDm0aTk3d6FpZUNbG03w/X7u9U6R7mhfLy3uLMyg8G+b4i0J/8fuQXBWjjV7tvmNH9Z6IWdrnV
rw+IV6F8heJkUYwQoM7CSQCwWQLLwxRDoZklnCPgOZC9K/qqtl3/5RZW6fktfk5LAbKerSEmubJA
bhrd8ZGkxX7LZfmyb0+sDE82uBXJOBt+XoRW+Md0uZllO8uj7qHHyDHuV2MS6R0bm2rNH0ugTwyK
0f0m6ujoZyV+/rjbAH4nWD364bogVfCTsOqnL7VrEOsOOpxdrrY/d+TWDEtf2gT/MtiIDl60LJ/2
/gmfmkiFW/vCyWyXI0ecTJ5v/2o2/MX7IjyUqtg9Yj0VnvfH5JoVSRS9mdxmiLUsFUub0JwF/XLT
J4/f5CoVcSFY25B0ONfrbASK5KfFe4tq4rn+eJ4qxZWAnYG4QFpUF5sgW21R39/U8a5TWb2XhpRs
XU+6NXpsCWkMwc0/sgZkj9Ur2IJkcIvuyrA0LtyZ2OR/iLvxLlWwEjxupwzNMmgSKTBLmsBGuwQg
nYVsX4hXEFhC1yRn4XLfMX/wObanTi3JfIcMW46c0KBnZfcE+edivvc646Pgfkg7Id290ydAoYWA
G0/QYHCE2ixDahAPvpnSUlysargeQkzIxhUqz84cKJkxma0GjKCLX2Be/uTX3JNn86ROk2gafZ94
7sNK7dS6QiJOWwHFFl28SNDkvfpRItNNPv+mfLIlA7aQ5kVK+BJgA5imDhFRF6vOShvEhtwuSgvf
r5bP/j4HRu1tYHRwR1P4CMsNq1p4pQmMWV+zXnabQWaGBEFGxJEpNMgx6TLUyXu2dm/RbU6F4Grz
X0JuwzGHzsWgNelqASqW9y+LDzhrTauF4O/W7QHa3G19Spjdh8sps+yD0O1zC6I85p/KiXqMa+ir
Im5M7GJOlw5bloVCUA7rcuLDVbAURc20txbtdOcEYBQMAPOLmc/Ulsp0e7FQF+fLVYzuWx4+7Lmd
F8ZcRpT9MNEVhVa7pDPOcYzD78/tQmUnJf7ouA/IFb6v9kzuJugq1VaAfN1Myha8bIYTy6uDsGxv
hr0yYlpdVow1wRNc54/TrP7BU++DHBNWd9A7vmlX/1YmEQhUveaD/uH7Aby3BLiAehvAifHl0FXt
ky/bGEyANX9PpA674/95ocsuWPxIhvTTAKeM1ft+x7ExBVaZvsfnQJEohYST8zNRoJPFwSDWf80X
PjSx/q5LbITxd/Qj9fZlvoK9Y4BhPakN5TovniqwRem0B564lwWqHpaK+F2kCCMGiNah021GN22E
f9BJXYwokg/zTi6nxfNTSSBOFSUpH2tP4UcWepDtOjAE3LBg+oCdkFx5583JTj0eOv125gZkCf7J
PcTTCCXpwBqPcFgBJtjyCrPHCj6H5nmiX6iDrxDd4rIdejfvjaPKgYYM2hZSRk3tEdEYx1MyODrh
pS+aLdVxzdaI7aekwAz3gSGew63ON4x4DH0RxlEOWFWFGvh7Bd+rQOEiBAR4U+1pEmRV3qGivDhG
lY+QHuk8pOyxhz1ENXSRbD2g07JP0SrzlC4+2WDrhsW1CGylXv4BNNGNICOKtzAhczhFP0PAw2Wy
nbAEI4ClU9i4RyiHyieF4wIO7cQRoOj6uTlXoYc7lDwgcwgHx990+GFBuMPgYVR8rSQZPF12/KHE
jtzAoGEt1C6a52byFLAGQbO3XEHGeDU403YUweq7bHc8RgdiGwCo4CuC1jc7mi3B3L3dwW3KQEFB
XHtVhzNn75WNvHP8bkFgUMXQrJQG3/q9y1p/OP24U/swh8S0e/p5qCdAtPrvwCymfdqrUJcnRFv5
pAXXutWxWPn8VN+6GtdefmN0X9Ie8qTAuT6ASGRZ4LhOrJ5kbbrQ+QXR9bf/+vdphjjM3zIqOSMy
3bE0RDnn1DVxyqq+ZxXqaNU60qz/oOT9rFFY/aY20v0pIzT+e+DzNqiuq3kEO9Cb2QVdvEs8obMv
mMP//Ma7nXZc18TmLbr6FsRkCjaF2d10h1DgUGbczjkNE0/uG+/zqqNeN4U4Q2mVYtJ1U64L+6CV
QJkQLcUaVI4qdsoSg9SHdYNtPdES1Q2ezNoOSe+jndndkWgEtIBPUg6vqJLq4894dkX0B8WGvwaU
iQCobL+mVpIvaF4ihIunxS9h9ajuNE/P1Wvhsts1JAKGbRPIeivBRaG9oAtjF1XT7sdLLobdXT+Q
Y/YeVLpWCXEyPkI/fgwRreQznoHee3ZfiBPhC3pCAms32XD7oeNuEsti/4BXFz4LwiL79GD9VnTZ
NqW0JqKU2P1IWWcF9zZHcO1OmR4IX/q1G8WnZF8Fi+fAfoOc1Jbk7hakGpTJczvcWAj6hrM7XHO0
Sx/7xGjMtIDyexOQM2JJ8jdkrjA3P04klbKGydk4F39pH1oCSxH2K5svRodH0ul0e4di7F6hgmPD
AK2fIvkE9TZwc9Uqsvmul2J/IvBCBQeeQY2wGsMLiwcV7qvk1OKSktK6ksUv5UTEieoBd72nBBC4
iijESraGbp1YBIJDHuuA9rwDF8DaM9Q1rh29llP8T72iUf0IOgfb2MavaOvIJaNe/TJZuRvDiVQb
9j/+gF5YtyJo1bB666Fa1RTUzSA8ELAutU5DZmvqTZZ2q53++0gysSrwdB53NsRGE6n89aCMZcZV
tH7S1z6Qj0tG4tRKiotL9G3pMBkvlW5vZHAz3zy2gRj9Dzsj0sxDulp+DaFBQgRzDyhv1MQ8zsNO
zx6Q8Ep4NBce744h2aZJ0EBBADBuIxqwjKm0Md+7aUOsr5Efweb+XckwSPzjdSoMjxfl13ihZLpV
0IyHcrZY1KLG32lqmqFOnD/sXKQ/ULkNg43GmGl6UJqqg0/rM0bBAL3+9vx1ghgQc30hHb5ZgtsA
u2139KZlSplSXY/UfAffmYortSGHNSiuIYghjt8cXPxdy7SdgYX60sEJEv8g29VkYvSCrShyM2R4
qrCdnnjKQelHJ94v+DBmfj2Yh75p6d2tgHxJKrPN2+ocsC9xWaYZnbxWORnK3HT0Ecw0zXZ9aGEj
kv6GV2JmZYBOt9Q47mgolgk6jzS3PrjajZ3N6hdZe677ytGitXEyolB2qSOKbRMkEsm0bYA2nJpF
zS2GFa/C0iLtz9MmX/9727xYat7ZG9pUfszA8DW7ORlmKBEpX7M8sLRFz/HFdUDiSVfO5nFnJsOe
DMTp5uoiWFaMVH5kR79bNG09CqYda8Y8NU7+dvYVfsWad6bkfXLOmUPKHglm6drmpvWD1DlRRshJ
M/o31C/ShuaNbFCFsbzPBDTo9N+8uRUDiT8XCaBj9+WKJQ0HiNw94CpqUND2A+1fytqc7qyLpysG
dHPuQFahte3k64p9rBUnUd9soKQnbNE93V2oravYQCLFpzOSmSPp4o2u4UgX8N+2qXuXRs5YTdK5
5/EyZaso7Xpbxx2DGQaCBTyhJMu8xshLZacytixLiTL8ReRLNdcJhVdOWH0odPOzZPUpZNy6uiaW
z/fmTPV86Cq5ZTg9M6tm3BFyOPmxAsZCNuA6NarDpRnKpwW7Zaq8iz5ic7q1l465yblX9PP2dPUA
FZq98IrfzxQ5D1ycKHHMY2S6ZetoMsrGqDVJ6pwaLDEos6Ig+R+YEvBtSkGxpOCXQW/DJB8tfuFV
6vK7m3/uE92/hz4AteWNyIjtgVdmi7ynI44GxYcSrSxDJaUrHSXr3YUHb91WaXL73kehyy97BtkH
6+rQANvei+fmhqnszcYzCruSA5zUpq/py0+6s1dtBt/N8y8T89mWmSb4yr5HpZiSycA1WiE3m7/1
IupxCh2bYIU8buBhGAdTFZfmBZ8b3dtf6UzNmbT46rRbHi9jZm7T4/it0+FlSt5TKvE3fBSJgqOZ
UR+HhgPQpIoa7zdAXvuUp/L/cYz1dpRU3PPddR1I+1xFW+8Gj6O98+6W8FKWtKeRnVPxxrUl02DQ
2lH4CynuWwXDVRLZC77/8D5Gok7YCKNXHKwG5G3Ymxg7f/QVxrJ54gL/98F2bP9M4Ro+HCzC6G52
/qHxhHJtujbYQgPwRzOxwc0s6io+vQxdRACJwK/lCdUImZhd7CuHU4wS5hwgVJmwWkFoSukOvGdD
d/Daqny59DcugaWWzFlkIK9EAMT3YeNR86IYq3FB/vMliEPHafGTpFSKSBYeSU2YY1Cr9WLyq3H+
dmLi9d+/VpUlJ9qgcnNVk33Jjx2bLZj16p0QbA6g4us35dFGG69L12K9e+oaAPWO2824wHTER558
I05R2Rm3u2FSoJxRZI+GKJq5qJYmbBWX0F8tQEYo6j/Mq7/zWX+pgPYBi69Bgz2ELNHVJbt7yM6t
bGcWDHYlXIfXI9gWD29/q6q+T08Vp+ASm18eCi0pwr8jWVPBMuGaGaH84JW1yeJ/JeQQ1JGWd5Yr
v+YDQvW0cR45iq2ajA8FvtOCOFH8XpdCrHI7VEnFmP+blDceQGZeJ6/6m704pLOSL2ov+mAdsKrz
C/3KMKGerPdXvNkKyPxeC4mJaHK1J+CcJ+2CPvsTnImJMTiYDbampUFW58MEExz6JZ5hNbpC+1Nz
jp4zLXEBKlocrqmYH7yPnrzS8sSkcBgGaoWssAABWCPbaHG5dKSNFmbT5UDjy8S+LooHy/nZS2X0
CDqKsp/8O6tyh9hU7BqIGG/u8c4/9DLJt7P15exbwt6Jmc0KBfZ8VsJNEutBR5fi7fTS0dEIQpK+
DrvZ7DHMSfCYCAYPpatUrRNctVx+wwnUmG/SmJyebicJMM+SXcWfZMkxDxR5MS8aG5xDDiV12LLa
hcClxRuYpaUTbsqL66MiZLGpDrgiD+1cR44kJBDavT85QosJK2PFitpnUc1V0q8ZY/0NgSeQYiPO
fkq4Kouf2oVJAYpDiw1gjmcj1uhRu/zX+SCZHb39RFMHj3LitVOWbbc2e9rX+bwuJ9dEIGt/qhwZ
vSyELdhKCJmQ/n4zEO1H+Zljx7SXlo1+pZK59gEZLELRaA7D8xQLbX3yNjCubGnPqvNCxsZ3JiIB
6CrRG0X9FlZUqSn4YZ4ILLjyYE35qVEvh/phpBC/JAK2Wr0Kkqgjepkj6HIBxZMdxu6uOE5tIrmK
bPMDvmLdKTVjIvMZnnxY/idSmn7LSUf1t5nmOrr6sR3MLwnWsESBOHMnUJgTZIEomtphD8ZMN/m5
iq2x/dgJRgW5rpO1cMFZvufYXyd/0QY+ry6GgqOdOCVRHdm04H87CPNDjsvcxtTC4EcVCATkMuB5
AmwE3mK75IOL+G4YsXSfwQ6A8iK/Dy+PuyZmt/eY+CoHakk3k9ro8ZcFpLK6cGL951Dx1NZLjkDX
bYX13M4blTQiTtFHC1D7wrcPjICrEb/+3GAKNT+FZfFLhhWDL4WbC8Mp5oIeB/uvRVLmjWWYVHIA
3thv8NxzjtmsZV9wc2zF7CE0IjgJHpRg9rS8YLXETbA3C0z4c9YQBFhvyrbltP4jtwaFkk+naVzc
RjZ1fqMOzJxxXi2iWQvDCbv4/BwT9cWCwmVk0U6MaJjO0eXXETlATU/JZyG/sSg+XX3AkN11MaMj
9UcJ7iDOvZt0rA0P54UKvv4kszvpoHOsaaul/HYB1VCgEaJfI5W75o3TOtlUndDbRKb2nDnNRzI/
2rHoQ9CoetsUEg1EaTxYLkfBkftqyALp024Z+ye6wqK+S2OLk0C5xV0TeWS89rs7zW/e7lJd6qpp
0rrTwHVF8Ipem+67ZuhV8XsTuNyI6KEk8O6SL02n5sWL4HKlIw6fDEf0eBh5XT4VTlFlQX+iLWV+
DyA3+tk9YzIR8nyAzgZWQDX3I0M7XKtxyj0xo0eWG208FiGQjmTtK9fVuPSUTJbJSJnvoR5U8rHp
dcVuwN/1mXxK/aV+LbN5tZ0qIZTvDlxIfSsRASPMVCt7afx5AJLZkec8s7VLsGdbJhCVb5H3fKV1
PgTrDVsRfClBgRieBA+p23Bvs20Ted5u3lD1VxbzkCpFXTy+BIvrQtzoe9ECMtQ55cfqtOheWfH/
wTMY17+meaXmhqGoYJlLBdKKnbJFP38b0fTwFxTb8sTv5CEBex7p8e/sxhCNQ0tUjfhaHasGBFEQ
aTcZpy6ZrgY0CHxlQS+bY/f1TzOWtgvywv9pQDdwU7lWg5OIZWk5ABYXVJ7ZUGMEScN9YnetVE7R
Zz/F2J/kMOrEy5XCIz1bLmF7HGgF9cyw+5dX8SvrA/zxoKONPBF34kUkWu8tMr9oYlc2h+xL44uL
f94fWvglIQYyn9+h5H6hDRUKq37bpXEhf12rW9lWjFZHTwp+XM7h8FU+07PaA9f3d5EeNt9a1ZSM
ibv9Mr71aOBs2uPVvWDr4e1MVXJ42djhzHVRdPgOxLA1kmCwEQy0QYWiYyCK2zg0swDNbpUWm6j7
vrSODC1Q4JdjQe2uaNWU6Or23p48DXi/1MTfFEhJLkWH6fT8WEAbg+Sazj52e5tka/1JVb4Qyqzq
fi4QHBCuotKw50d1fo3Hr9xzSVF89TFlcQB8izX/HPH8XSEx0s1TBZI+qsitnvf7uzPKnzozC+2d
6acSwQXwgUXpJ3rrJ6kIdW9uytHArIZ7WxZyWAMcD2llWDRxTYsv1THxmj9b76fF4WRs2VXp79fm
TUWrxy3Y/EhML+2xW6Pt8y38g8tf6hzaRiOw3SIJqUBFKzXdzZI3z+SgDzG806U6xEOSQ/BcgH2K
gablP2Kv0Or4N4xWXirg9J1k+xy5hmVEumk1BzgTQ97CKmM7U5M/TfWk2OwBiQiChljWDX6YYP3N
oPCB0/LxEq18CvPjfJhQdzHFopKXkxfvfqHjIOoPY3PW3n2cy4I4KfINdTiM39kz+RtizJ8XHOek
gXL9eRktO5sVE67bySW74OW2745Vm14m9LjnhxWW/h2Pnq94c6hVp/YQeEI7ALPT58LL7Ps7Gywd
/ZIcpRZAlNLUyjC8Bcww14h1wk7Skud/suEVNm7FTxXPpUkJ/KVYCebKiMb4UWuvzbh1L4PM9UWj
GAqS/cpd5yzU09uJCohPvDmxrL5j/TpyNbpRlfjCH7r/NCSFLVQxfo3GXmrE54rlKYGoa0Gz2CoB
v33Joy8Is88/8ZyYZ1Z47QVQW7MIHfjUtUiispDYXQU4GK0+qbnH5/MSa21PuD3Fd/DVdwrekJ+a
YkxDSXmsfEFWVNFQIogXoUkgaVGfV11Gi4mzL5K/bLTII15JvKjDZgDaFVpGjs1T9UoN5jRKw0uz
MzzxTWId16uwfFj0NwZWZfsd+v+rDPidze6dzOWDudB3UeQgJFwZfNCP4JWQXmDx/EgB4fSg6TXT
Kz3bw0oQ4YKL3k4QZlqZA362bNVSq8JkItP45JAzoxpxCdEyZODhciwuDqr0Lq8BkQPCntdvHVqg
bKk5BTGjG+fPc8e+CImuKXPVwYQG+8iVZvHvRMqBCCGa2KWsRUZu0NDCKQp7UD3EzFzgkfYBHijl
sQr1w4X0+SLsQGLreHPKjqJNCv2Fwj7CfZQVTvXctuoF45LVqS6g/TFPwRymRbqsC0USefchHH1G
nwaqYY1YNECxRCnROYfuQ0eM9hM1KaluLKLIqAGEx/5r/xpBYhijlcmUc8q7bGKZbkj4z9c5IDSL
4jo/9ql5svMlgyJUS14q9g6MSU3nDm9rQLIj9stijmUHNAQH0TDjwgenIlcUUSa4+70vaFg8EQg7
MshD0zUovNUKWYvXqw7WpkuezyoXo4EyjPPr9p7BglbeqoRbQ26wYcdkKgLrN/LjIVhFcQf4fnBD
2mkiKJaEYFpTJ5ExzYv+OGxvusUdfsZy4py//f16tPgS2RxNdvMuPONX0PjkK4npZ8plspzJXD1u
aq2DgF6iGytlfeAcLcan/Q3qLuExYZZMuW0OraXx65jt+lXPQe6oW7PWZNdqHzBxsPy2teuOjHNL
pGjeUiZamGkOgT4h6LEyrVHcqOwu8SP90FvvRXXKoemr4Iomy4y+HLyO/dHCgzjxprEAyfgJLSCF
+1Jlhckkyi2EYna96J3WT8oTT4fOERr4TM39TvSy6ukeqix0nAh4vxGPTcCBLGB+fA1M7lrMzp24
sC2AzrMDhbCLXYl0Imu5tPibo5GUTJ2+zJ966v/Jof6j18xHEkrYf7O/76wb4d8VihjZ8jN4a5l4
/TaKbXc/0aE6KhQ+UHygYdZipEuwsOYqEHWHFj3XKhiQFWozf9nbeeXYdiLf10elMCxXKi0SgztR
BhWUeo70jx0PME20dIlXu19K2ndhzCXBXAMFlZgFKIswNzxWAtOmiv715OKAXpPz1mGIEtqwcRsA
WOKkfvBK1EO8U7l34RuC5Hfz7wAvsEuk7tOJGL9eJGoueHMV/cOCN19xhMoaejdsP/AEnw0usc2a
D+Al23WTQFDmEckcgeoyTwnXjXGsB5hw812EGREHszsRAfuX/WF/y6bHBCzW2LLrCbpQd/YKu5TH
IoYMPqzae2TD0YDZwWnB6fRnsOV9syiLzqZJviu7r9XdTRIt0t6sUvh9DDEFqmwTymr4YrWjienS
Mk6uLSqBniWHflHstShUfVUlWfTcXy+9d6povauZd8KdeQA5Hz8gSp1nefCqnSrG+IVufeyoaArn
MDpuvBRJVzn76pJGuBKkjsCGJ4kLWHKTAdfBpR/4JlDbnqCaDnmVWUyvTb+7knkdHBddTiYZDsjx
ku8+v63la+9nsAYulB2u9O3VL2XMnTSK1Ji1XvaliXzeG44zghi+y0NsPpzhMrHayxfJaicpNt6K
fFleyY9mJ3ZIme5Q2F1XZ2ikf9jUWAcXopItzMTJe/Hl4Y19xFTvzMC93mYfzVPkw2irTAl1N+r5
vKbm436VBLejR7QUuO1N//ESzLUqcs2X7g/rEkcLoK8O5dQl2yiy252S0+K8xEZgx+4MWMEEWpT2
vo+u9FHkZcvwKMfIylWbQSXaJHoWcAOkJnSQDOou+f43NbBMIf2rL14/UZbY18pqZfhh++jgvKJw
B3XcFzd7zmgdHnEgdPjDXL0f4DJ0D6He96ni6nCEG3luFMwK2m5dLTm+scXiAJBDUd2h1dd70Xdg
y3gScJjUeg56faZEz2UGPU17j1grcAl8cMICtui8CN/KbTQBGHVqWfCvt/7dtoXMGdJefk8ptWg8
zcjEkdi0Yr84TvTh4Kxrcg+scdkViAbgqEJppZX3T9AaTvl0168oOoMU1sLoZeRBOAQQe9x9Bm7R
y9tzQacRrtbfx2dNiiG1/QodBRvHddPyGAZe8qY6YKHjTeQ2v3RJMF2PqszBpqskIGmmYh1i+AP4
XGOY9zoAetl+gfRkdcVLJvxIwivGDlyddqidb7vDuEq+QaC+p2L6r7ws77kyXOcR/rbOvliv5v+O
vZsZlbD05uvqvXyi0FE5Pd+196h6orPSyOO6qrho0Ozin/9qGDtEynvL8K4fyu4RUmFOji57S763
aj8I2GNfhtQIvXcarF/uWxEzvOqaiolZj7vT2/+nHY2D0ASXDwapo5Nmc1emmOsMkNon8xOZPjC0
ZCJByedFr0dWcnqQRy9KGePne/h2kdACw6xf4LAu3rRTpzP8Suga9PxIkXhiXdoNe/sajJeSWDRI
0hOWCsInXkzdSCurz5mpx+W1mnToV0KXEaWLHgjzh9d6phKLFmKZjQzIRFzBkLCj56Fe0MtSH0ag
pbnMPVAjLGtBcCg7n/ul4XfrvuaNaVfOO8EinkIkvzD6XMaD4XkO2nRy/7mOwhWm1YmsYtVQpil0
/x3fMNaD44hdDNlUudjSPl7QEgDL0QB0fB53ExL4nprlxFDxQCeAGo+bcjbYt7XVnaOAE0HvJnGw
LdigIYtTkoHDDanKhz9XvUHk3fYurAnNH/yqjgCy3346eNNYh+K21RJ9m/JcxbaPYQm6POIwR0Xp
x8+S/llU3wNwAlZAhImpQ4jeMmYfKVmBUzdPyFSGfm3HrD3piYCUPuGvlwCfFp9UZ0zPfi/D4xM2
z492Oylw0LsSuPLv4AB3C1aeqy19jbRiJQ4gnTx20KIc2bbUFSKdP2egOGHAy4mgDWIdYPyVS75k
GAdYGD6NT/GyCV+8X+VTGQ4lZAAh8zOwIKRPN49M8pP53DN8328qFawShS3U9J/VGqDIsG6AvFrC
6Ji06pebp8dgmqjiTQ987khRaWUbnioF4QKKF9sdbEu/kqPonWLZue1eY8MvIVlg4H6Uk4foUIUl
fGVhhjezkdKD8TBIQd9jxd+sG7Uc67Ns+TeEtG64+lmHSGloVkXcsiVJGWI5oQWQMlWJ/eFVLdOc
NfboICjp1AkJngZ6JxfvVnkaFkvGaOGHqsbMSX1Rgw8v+lQCKbIGIwknDPhru0ajahgXZElUmFM5
zv25V72RFuLj3yOLjVHrmzHwoDcvKHwEKlxa5y1b0NPdK1u9/j1p2n0/7DL7k7PYTgL+jN9vYXJw
s+5y1+kX+mSXbWSRrmyqB95k8MOmw64SBbPukyocxMcIiGe0ePGp9lgwn89/lWpUF9cwncBqPoOn
s42CNZEsNH4yseYIQqnIAwk0GTv4j1cPeku+71JytkLNMHywyETxjH8IJIGjFtPqLFIiTVWQP2QW
6BFelY5G46Nz0Mxr8N0ME3+tc6BJbcTmjNp85VTSZHD7ccDG05eR4sBqX4RoxVQruDhtoieMMJQX
Wu1/1rn3zdvb6R9J6dj21uZoUZzKZz/mRqVfhOxwiWcS+YhTiYFd+fa0EnJrtvF0ItUEbxy7vwX9
IN1iLrGljRm5eg+jPsLuoxNa/DLaf4wXiqoJql1tESIKpU6ksN8orbbxGEnmmK4c67NNZcU4nR4F
gPQ0e+PFn53gRVdDpk4UY2Tk9pjF4TzfyeTorXMBEQbyJG8PTkG2rYvfCoD6ME4PafnsyFG1xYfl
vjGbnOTaJ+VFyAFpNqD8TpYZgwpmO9cyyJRUJNNpip05TmUJEIjBzpsywSRGYuwEMwGHXrv1Vbc6
cVdNij4W6JglSXvHysHvWPawDVd7fEnWTUS+d3GFFg+iD2OqpRaZI/ApUJ+hGkVBsm4NmNmylBb0
PDODFszsB+cV4ZgisRP01HtEHMx4vq1AVuouyxQYCUCS7y8oernmuwHxGhWdFdUT71+nK9hgkIP5
WC85Q9R2ZZK9z1bdmr9TSTf+TEY2zDVJCy7r+hLkF36qW3xtKmfbTmVA9mnphUAccKDqPjNrGq7A
DfpaM8y6siGG/OYP0LMrk+icfqikdP1LqHb7JK6m2Sz7GEevXeH/uls1rS6Jser/5Z7THnPvdFcb
zZY7+laYPdfos0k0dI8GIZUFumzHJOZip5WyeUKgrUJWlcBtE24+HuQtPalx+FffpZ5xruuMwb2w
jj8kOGRZMa9a9XlnR11VZjR5yygc2Nruqg9YQ1AGy2cf9kR+Fh8da6J0md3SZWFZFt3Ccu/k7JOV
DXOHxxhqIlQHyuCz+6rB2L674Joao5v0lrppAJnqxhd7VMeCAxyiC5oXPxqp/pDHd8gcWT6ABizw
nLQDm7rqskvFfbGHHIl3rAQQMUWE1zvWBPK5bKtY7JE/lWe9TN4QqDCKNs0momwoZTq/sHMU+Wg8
7WURblthVLeJ24D8clZyz5wMlFzX+ztaBTHwAEvXXNq+jom4wWxt9fW97hbAzA2omn9Kp6LHZilG
E5phtqGknX1I55tt6Z81V6pe7c2e3fbLu6IlCTsIylfnUu/JsiOm891qlilQT66keYV5Wgu7tr/e
TpIgIKIH7xYBTGm7sGahcomXWsE19qu0RUmSzao79XEF2W4k0n7RzdIxjvtzUu/Ct3EGeGB80m4D
bNbwWxj/t4ASCF9ffjEKfWa7dQ5I7a7GUwl+Il6COtXm5/R4SLRTDSU7HxNHHUs0F0kPMA3t5Knf
YzJhceOd5a5aFO/CH6k4XP4dK4BTNnK81/YKLAX7Gv65g0T5wsj2e6dH150v1uiodO8/nRbkk0Wz
1iCskZsEwr+1j7YCUjWO3pc8jXDYgfbxetGXGPpy/JHff4b+nQKk6/Zt0UNbEk0Xb18r8uaJrG6g
mNqWIUEgrQ+em2kTv8VtmoGC8PBvkM/lSnWTfgyMjFo0ANLm6wdQnYiRHYXTmNIClGHqxzJ5x0BM
UuwkciaGGtjLqmTY78ELexcKBFv7Mh4WqU3G3WJWu3VQ4Hnsmf5WYGNh7DoaqAz+wtwzmzJZt5bk
j9U2CnTJIrlaItgOWUP2RpSU4DLiF46N8XYuQQb3TtwjrhHeIwQeajuJXQ+/PqBNbkelI1YQVIRg
Z/18JjLfDN6+QTtEvUK9B8eyjtHy5Atn60eAviKrE6BEzTwGvxCMJcZ+gk98C6plY4AgzaXw5qQY
+apF/8NsRVGBLOe/ahDgdot+GvvHlp+RQeeQSgp8DzLgRxbTRugUlxC3iXKQto3TZlW/lz1o/r0x
Ey7ku3+w4z4OG1LznnMp82HQGq6TDd89Pt7AS8u/1pnTOLByhgw3dcfd5bi0U7awuDHA4Iqi2OKj
9oMwvz5WPQeQD6YKwRCyo4E4VsniZ8W9w1izza+YJ9+hEXg2qbu+uf1c7lGNtB4S7qWaOnrXgTE9
CkQA9XDy/B5KmdfiVWZZGiOx8oot9gzJHXPN8JKB4lk0QPcnoiZEziCauHXMpeiMLDwKEDBlOK+c
ZhW+9PTafeB5K/yQwU41vYCM3o8HAXl2Os9DNUSxkAw1SLaIMKrBjEseIG43/BlfzlhI001B6z2m
vEPOXsn9i7ykwAf32/mqCvF10r7yVsc9GIjW048pDeK8Ku9tUov87AhZg94Y5lqzVNFm/2UQg1M2
rp8Qx+EMFbpXWpnp41fYfFy+xwXYf2s1tVKgGtGfnA25Dasyc5sQx/pNBeziAXgQrJLAAaeSQFxl
9YeSh54nL8mNDFW82l6HumDCyyXHXhTVpJBVkHcpFHB2QPvNNK/NyFMP9yw+44FaTThcTRIE+Zkl
rYeyJpD/7U7ToofS8hMLYufDpmLdESygwHfr9ojIRU8m8l2LjsvoAMGsBluQtUdrj7WSupKv8cPY
aRWtZ5KtP5t4/7CGMZxneFdGMSox9csOEjTx4gz/zFFMVww/D9LLaK9xZI+ddpZL5g+e4eAi9XUA
SrH87Be6dqfbxYsoUUYw7ga4XX+g9onRoXmQnOmVx9iEkrFFhabfCHlmIsg0aW02ShqGViI8Xim5
ENJok3/lcWzwABdPkkEZ2i3UJsA4XGpbX3bKv8RX0bTiJGKPhopmwaz2cVheaalOFTYxAX4CMmJm
/iM0cwHbEM8zRdcaJGjzupKHAc2yJyIN3fjM8WYgwyd3vFR8QswyzkG2tf/bwXwR+x8jlO4hEMUP
3RkVUB5UWAQp9HruhFGFr+QRsYP9keerpUfz5NHFIM/3YdccMao99Gm3dqOEMghioPFKvnuP7K8Z
Pr+M7VCKJRQ8uvWZrM+w9mx7KDlDCnKHiDt9goiagjUXak08r5e4UF22WtJRDDyeTVCyvEfywCUv
eubmsqPu7vzM1q7yy6EF1V0qk6Gp3iVi9d9tVuzfn+gY72+nB087VgaTGLpH+Bi0STEOin0FJBjN
Vk//svBn7hw392kOhVlsBGt8iVWIsc7tlvODxLW8fJlLU/bRdJakiVFuTV012nzKNZIEZhmUUV13
dvpqyOMs7xMq3jkbv6RJS+qECrGPlzRzXXzWIl8gfljU8lsrZJ0wwN7Pe13oCitMnk7SGlP23flK
MO0Z/cMw0B0hFyQv9e9xOiL9Orv0J3hHIdECPJh5cg7pDR07AUa5d+iF/LScZh1HH4J0KhEvOh2h
+CWBInzCNpCHdI8UPEt4Wm0+Dao2XW9+vQ460cQpCy7PH47kV+3AJPFJOUF/7I3/kcSlr+ycctLE
Y0WtA9XZ68M9NDsVVaIRse/reT66dAmh5aZkXfY3FOO/gTUs1+Lqj2dDGwdvvJnCO/SnbXikbPBA
dJMwJgt93QsMzh5Lo3LJAIlmCKry/i7T0+NuJKMv5VRtFx+x9110dam1ROERrN6+spwWO84vsfKH
7iOzC3Zm98sWmUwkHKBT+zMsbWG3W05p2WuINs4XGUu+3myV09Unt8gU1JCC0iuDasZHsU3iR+Yc
5ovTrM2k2oKoCe0lVJTpILAtYeASuP0h/GHvOArdYmdRjgbLSSgLJdjDuRcmpZJjKo3iX2RNvRSs
5xsu846Nc12NNQ3c1wP77A4g/ZC5D1nqO8FA+Z6/ALBZwEz3iZKSOFt2EJyYDn9yUH/U2jjlLn0c
GYIJg6uuwfGJkYFQIO9rdtVSCfj69Y5bIFvVLOW+sj0GfIsYwfDqUoselCfuFHoi570sTmO/aPkj
QNar/HgBMAK25gFV8zaZJzVGV6+3hJEa68SIBJAsIoFwl+jVpphtxHyGA+HaweZQRJc3uOKTzsPc
422plHA3LhsDDm98Mca84KLW7Sr0Cn759DDbBknnwjZOYxSmt+JGlKNHolNOlSc5ztvl40qkQpde
/lJMnY6YEpTsifA+30woaNbtz3+4I8iIUoaYdyp4b95bMCodgnEd2YPWL8U2xJZrTP0QrMBQii75
PKQuUrfRqofayiphgbJEOGrfSgTBKOv/u1F88ead1PqJEangm0MSdv7utTERo6xcxIQvqN01wOa3
7+jUC7xpeEg2gJPUPNMg3wgV1Jc9+BjdWHKoE6c7DBhCe/iCvYtVJGWsn7wYTS3ujOTPWlSNrUX0
I0kL8ZmAYw+3rd7j0aOS9/F2DOusEHJBm0VmFGrqUBukEFbCORRibn8zTQCL6usEBcGlA3/Z4gDB
DXQU3HVErTspLpYSwLRUemxzUQvQ4Jq38yrlSUNB+TslTMAKGvOKbfL+dgGJxNx8Vm9FyHw7kmc+
PlDrhnaA7PyDmSA6GkmfrhSgTHA7Y4LIcKVb2qph3Q9bmPSfm3zaJruP7c5X/lPxiy2b+l3pFJrF
vLP6q8Q81HBZnXF1PG87qgE/eBM65Uybvx37LlZ1bxZ7B+rTtCh5C4yEE0aDGT7N5OZwemg2yP/K
ZiNqQmAkvQNrmnyMQnj/lFA5pIaI31lotQvwShbWadZ7JimtSQdUYZ9JRSMPrHGUz1ALta6PMEUJ
TNHp5Mn/yHzS/J1J6paEn1hmMUFRf7AFROhh4v55dCqIlaq7bZTrhAdEPhaCsUApzARniXKoYNg7
WLmuxfBvzt1AVugLJ5LRbMD9w4j+D2uxkO+JK7vB8oj3kusmOk3N8bUf3gAGsSemqHFeHWwH8Tyu
90cWImCz4lKse/uhXM82LSuW5eA7+Y/bMTkAKvEhNZCLGso4jom4yCiznAlGm7pDezzt7i0myH2a
1kcGmleYbBtuknT11TWp4aDHyWpoRExxJXd4bW9vMBXiAZvpPuJidZl4dFMI456sD35GIId7gPGV
7ZlVo/xEDj87vFej8A0DpJ+HHaf9rygFWZKr5OWioTbudjAwSZUBCpl9hDcMBdB1AYxHwC8+vPkH
7pzZWklJsuu+cP+rwfNQljFDREKhhsFsq5WLQxLkT2HCe/vkIuAD8XfplTHSymJ6XG06kx6EyafX
qKl0VIm3SciBlJDikPs5ATKQdtTedanDX9ysdLnDgxcNJnOKSD3fUnt94Edbul1qjYFbxMxUUi78
hznjdltYtAD/lzHqj8YZwAx7MsAc85sHRlK1a3HwcP1ak2EiubWx1dt4fTXVZt/fJaxnCZAKAUJB
SDUeHD7WKAnsyXgUKGKy9V9ejkJB5ezdAUhmu4hNrvMnsanO4a0o3yoa+h9/hMc9SmFfSCObyitI
ZKh3kL6RfB2GbsCo45X3Ky4D1TuOPLa+RjP13qjD6aQJBdpDoA178Fptaywd2vyeLN+fmBpfQaQR
saUcvO3PpgpJcGwhk8VeU/dVYoU17hhqPlS/poOjIS14NYzc6mD8C1pLLzddLNtHP8d8PizrXwFm
aViUc4VKrV0ioepvYte2RQpZYkVdA+VvbvPH4/Z27C/KhJjqXopmB8/6PvHEaC4BZIRFI05yU7HH
rpKeVQVEqn0tiOI4YmeunVCfyWM9FsEPoVa/+I2pozpa0uvuud1WewVMHOmJliFCcuTguL4tlGaf
+BtLKq6W1gbKgy22QzjZN8E8KeJxpag7lBLPMUUYZtCQECQGoLyq6kTB/N/D83js/+Igb08e0AKH
jE94H/Cpch/PGlijkuHBDmMipc/o3rPcuwKFvTDnaKWGMN83K1dBGnkiaYhV/fEDb+6T9Cu7d3Tk
S/zuJFJiOg/bWel0V4xsWOfLbJmHht2E384GgbWRKzQwPaNdCLWxZcUUS4nudLnWl0hsZ6HZK8u5
6v1t1+BgrXUbQxN4bFSzLfrsP0l456cvQzy8V7n8DN5zy6r46eKjxQKLfcLlW6qybbDRF3qSrUax
giGq+8iIwAK7KravSl4b0GZylwL5TbjIPKSmA6kPKt6pvaTL9KaExdXRN1vHAIqSHvQ7acVU2Zmu
woY6iCLo5ZKw+IjPH5CCWcj5pjBVfUqwUtvCFAWNn1mYpd0IfUdMJLvm7aOcbxzrXT0yhXdyHpar
ZW1DbrbHoyU0ISLDBK7mjpsB2QyiBPXiU7iAcald/O2+hej5dk9R+abk80Hjob16jJ67xGvJahNv
hQaygJrJKAiQdoFeLSV/ww1rVj/hCGaHg3682nDT6NLdeUKAWl5h0SwymYD2BGOYeuIJCbY41YMu
fS4AvKDQLJfWdKvg+aiNyVlDEJJQIDZRxhu342WqTUdwYdSiZxVygdwxHAZeBG1o7/nMg0E4XEy/
FqG7xCIgjhAlw+sfZ4l5pQaRTLHLPNmZs3kmbBhfE/NpEynrZx0cegDD1yViO5oS/pBw4wwOdaiY
CXSLVF0ap9waCv5ShIscUwQeFwQByyli462kiPxCnY0sSYOc1orExkeFsxHmIjzzg6C+Th6fWsiv
4EahzLeFN000IqP6SQ7oK6VQHnwHeaga6HMfs9QZ7cUvmETODx1YFCpZ6G8Bw67jcko9wrBbDTrx
t5oCJifW7XpWAIGQq8NZlDThWFf410tUCSqj3aQsg+RlQVXPfGazDhwmYxeNfXezKQ15kyleoTRS
gisSEpbA3Ft6JmeBumu64FoAr8z+Qcp1BRCbiIBhi1QN3kN64l0pET+HixzGixptpbRqcKdSUbBU
rOmiQFOGwlPC6fs+CaJZKdUiv/9CXfkoXRDsxay6fDqe0K02a5HinWZoiLQqZf/vTJV4RO8OQhbT
oGNwajDSrsMJqWnu+QRC95yGzZB7CpNqmlBjKhOc22/CLPOzzEw3xnJK1Vsrs6QmhHm+jAHtf/1z
aJ/y47MsoECCJTttVFwJWiWmHxBBQFgWcjWb9MAwvNaAwz5f92zi26jAFeCeoSVBV6L/CnforcFr
iQKZvJ78TwU1jyvotV3sFgdcqUV9LBu4AI+YK8aYAWOZUgVGTlm/uc0LCY1qpI5tSzzKQTVh7kSE
/NfaIYQg/d4XwBjJeDGGdqW0DFguOuupsY729Xysj1h1yxFs88HDXLrZU6Yw7V1iajzAFED2Xo4q
Sv67Ss8JAnejwJM4J3OPzGb1gTG2gllLFNyvZWxUdmvxABbK8/Y2ogy078Egu8Jxz1ogdn9NGdGL
sTYdTZKzfrvRs7wSduim7HiRZz+lifC91CbmxuJMawo3u8vXgnB4SRl7OBBz9+9qq151IQCJu/1Z
5I1Ho0fh7IGWzwc4BcqzidMwVB1bpiLUy9B0k5GtF7y0CyMYCiOFwRXj0QC5faEi6mzP7eawpXsQ
yZ9Evd0tlDGLmx5TrB7qrYMf0G5tRyaabzHpmdliB4C1NHBdRkN6pUZSIBASf3QLGAEPY3yyHu9n
YObaBKZ6h7fcQ01j1v7zuKXLZMj9PInvo2fY+YVbEx9I+L81I98zzjx7/uHh9cAcPq/ujuEK9+3S
vknmwNT3QwSLmxKpZr4DIoJURIjySxurRNOl7G2pl7dTZFTDspsJiODB9/gjqP/KPHfmmMR1bOV6
JmKhP0yH8k8pJy2njfQNniZpkyfgl2zxUwieuUqUlrxgmogi/69gVcTNSRs72lKPRppUs3LqkvGy
3pE574NYYFLwx/wt8GG+WZpmSMtG+Khc8pcyEZpngJYg3n7yBj5SIG0FSNWtIePqCwoTsBhbeMwC
dp6JC1FL/QgxOLEij3y3ZNMxfBsf5mRRcT7m5BGOi/VwyZhf/T8ohuQgJJSZQQP2vhUt5ob9cCVt
U/hKLlgLLLXje2/UPEUNb37ILOAeuqkY83hb//PaB+TMjMeTjcynAhbhYOiKPYUjTiuBA9/HbToT
Nrom2LzHxWZfuDssvDMQp/KRQsw9Hf8fxyXuHnIPHUpqwZWJ4skGB3qwpwHJcyo9NB1XseCQJxzN
O0zECeTWKMZ9urkQz6UXrfDNg8A2xc4snMethxsoB8RMKS4tr+ivyuVSlU9nJ2Mkf7FuUB+DnTaz
y6DBTCtP49FxiWeGUnWQhBbsFh9cQBv+VJFpFNrZvQAlVuOCXv6IBM4++a2UdK9duQUDCk5a35Gp
p2cT3VpmOHVdjvDW+noGbUYr3nelDnVkNuv22deAxwuuTfay6tbp9iNN+D3pr1ZZPKzECc2/dKc1
qAh9kJN84j8C3mUcBi2egpHZ/7CqyKMKhzbyTB2MfKXdtzZ3mFdM5w3oDm2K76yUpZFL2Uelcw7A
is38lXFoSj/F1cf3T6IfTPWitBe41eTc5bI+CNETCRwGs+Uzksh8h/ur0m8JYmpv2s9OhAwQbj/9
5jMBp+5VEuJS4Wd1byPeCzER2sZNUU2Qco46aGY4NElV96TrFa5NbUaIpTXIof2EcL7WobpXL2eC
hk4p5LQgwttnbAJno2ste4aPAATCSI4VkdNvEj2b9V3LB66nJtYJwzG+CZ69ZNcg271u4W/e8dqk
GmR8cbThWXEK3KL1MxPN8nv/acFGHXAPa0LB6kTFZLAKCYwOgGX8x5ibH/C20TrhTNIeeVzN10nL
zLLNNZl1bhU31oeBIkuOwF6PmOD2S0YGsayFaSpOVhleYfOT+CvmXlsf5XZnFHuKnCC1GWbsiPri
UzAutwTOH2pDLb/JtpGfj/eBEEIhf8T6XFCVgmZIY/RrohOVTtCjMVIkCLLtH17CAW1Khh1FnMFz
IZ08q8fFifap6gLAXFeH5tiAFqlTTnSgnaBy4XazjaT47DRA8x/wzpGtSuVQz8pyD2zFaE1wGABU
94uVxXfnxCINv/jbjftvwQUDHN6ZNmgWaNbtVdD8hPat2wNrPyqFPYz1A/RvCUQOhuvRnqMdDA2X
p7riv/E5IJx5pOanDq6LZ27FwAECLV4iF53lH9wLPKHYRXNM2VU/rhge2eAyCszC/R8KiEFxbkKe
4eL5ktynJZfmZAA0ABLQtpyJRO4+Qkk9OwwyaV99Tnm7HPlXzX4vjqtVEdUbfvQ2Xu4bHrhw6P9i
OQTWeAJlMk3nlrb2iyhPcb/XQNZbbDeacY+Emo/v79d6208JK3dcblUYiHVUDNNCPM/E0ClOcw8m
KcYhyI3/6276PWFTpS60Gwm6THVv1MhYOT5tWgmeJITaImV7DA4fOjBC7lRt19hhXKVKSp9bt5D/
7sh2jaYVOdkib7k45ZfvN9MjEtXNy/sJcVDfVjPdMUd2/3CQ0cripP5KZI6+b7crMA/AHHsF12Mz
D3ZBClVGU0n6KfNADDJcZCuSo/Mo0S0QpoRn8j7ek7+pXAoqT+W4t+XvKQPV1wcHr6lk+8ixhoVA
hrmtGnPjsjFKvc659+g/UcS1/YGvgX0D1ZdbtGFtHiCn8cujLNCI8nzRVGlp0W3wtXyIPo0nLogq
IbbQsdi69iEY6wAMkiIzjsYKjk/iOj8DMAYYrY6qusBFP+r3TEOUvyIwHbzJ35cXEIhW4Wev6OV9
Mu/J7xGPH000oPbvI/146p4DeGqUmlEAtFRBPky3cNuiHsL13ePUEnm5GUOQ0Fr6yTVeKBoHPjEF
gLPHoGRbfwLs9MjXuIl6lo+Rv0AXn0E7pNAbjBajlo+WezqFOFIeXtg3lLA99JotMtZc3Y7Ibizx
g7ByUjJ0ANB6GeBzrPOH+FJ8aco+9Qh4Ny4Pj490CwpJCVmkcIA6JDSiVg4XVEtytjKzMteEiO6Q
Sg5lt9Q9KCuuQbp/iC4jF8C5o/KGoVrciE6tjKR9HG3jDniBs12agaewLVwnD5kFRIFQ0ftkRuZI
g74Tu14O+6niMC4WIRUzIK/mJNVK5Pgr0dfdW7tfQwC0MNSGAGGvYMLPOd2SmABy6++WVOML44ng
2FvtCZx3dxW9svrWGAICJ2FBi9alfsnECj9srnXflI9ifpAJ03PhLdN7ITujX9E18Tu+7KjDULDB
7kwSKtrDVOMfuu3Tu5Hpp/IbmB0xltQ3Xd0NXD03qDaEyEQ/e7arbc5VPMTynGSb2M2LQCjMkLjj
hB5JCiFi1l9QfVNOBPfvAWgE8byi/wZc7DAu27o0qAp5XajSsSRSta6dYawCiVmoho6symL3cimL
BtnVcRjJoY76oZhDiDljqO4iy9zAiDsDTWRb7EDokhxoXa7ueoqD/QIr1e9KOXv2DPvjDVRqYS2D
bJx+7ieTij9/17p2E4LDXWL+Jj8IDVd39LUHZwwteuPQX1/d0aqe5g8s36bNQto/pofTjgoVZ79m
eTa0C5sJntvYRChekhf2QG9nc+Q9oxd98GVUPa2NXSsu7Nh8hm8I87n4xhYmLWjpD4XofbLM90bu
NVUIwqzS3nmQMynV3MouR0OFM/4ORinPvRLpOWJ1/Jofxw1BI5fxK4CnnnKcnQWJwl+2ENy0bieT
v3I9OTRCfJz46RJJYDpFHLfAN0yMb2MFVf9p2W+WjDL6Ym81QSng4+y5wLl+3VxHDY+YuHIjrLw+
MaBAENw9JRvXFgqygtiOYDgTtD7ugQ56Bw75SqsNP2XBsed8Ef+W1GyihduXeDrD5EBXgrQ2Nk76
hsar1BEEEBlChCOJdplhc8LsVmi7Nujpj40Q3hgUu225HsmICIRB3AWnt9dH3lnMBJ8Es9bxujNo
1pyaCuCwm5rbcah4jyK4+T9Y6e+SHj0bj3j2OH1HINhKKB2asVPdrW1aZE5IILkFoscH+ys0XApT
+8Zs6o+DbuSe0o5bfurizBUQaegKK1yhuTJfVqXxn2mgG+4EvUz+p1yaxB1fzXCE+H7BHyobDfkf
4H0Yj+6VHwjhP+8U55fss5FeDnQhMY3XPKSjQ8taKULfte1fiKSU60yJgkDHMd7QGHJx10ksW9rR
EaEhXgPpTQkLOaRUISTNy2rfrfs4tuSRZCHexPnyj+zYuTcuZQ/vIE8QTQZTVgWcTyysFaJErdDP
+i0VJ2K9MHVNTRfKAW1+2+3DN0sXZvs8CVcaivXaBjZEM5cYnoF+LEmvqzvdAOLwGDb1DMxrbMYE
6VshCiHpsa4njvtOz/j2U4ouXKJw8w6xEinX0vDNj6Yj4LQnUtDB7LPY/dRVy+BLLUV7XIwTEBob
uae1tpvjOiEJvdcj+WCnfxfBz1jnVqDCj/Q3s7beBRjRLR0wePrRFr6dtCuqPo9hE5z6ovRmmmU+
9xgettuo8q4S3cMb2lO6namJibQ2JWfBI0TfIRBH+SBaypF3UHCKbxgH6wBl2aodX7gPPTOs1hNp
oAaJPu0CoZXJJp0aHob2PoUzEDJuY2+RR3D52ZXVwFqePqla+B1m0Pz3Jl++ose3/a0LvdZPgtez
4Iy05meMnbcdhczN3nYDIATe2KEahVTt+uMwBcDaUEJsGq5AWL9HHcsK7wzccLN8/+BG2EwCdPLo
D6h+SqPaT8q5YyEldoCmeGxu16OZhzetWiTJ1cJONo20Vu7CM1kWFN7xvDck3VxRupTx1bJCpqAm
q8IT1Pg2K37fcthXokQ0AR+73bFMWXt9qQ8dr4Fqv/Z0slnj9rVwUeBUtQyUcVA3yKJfhzVBqWUq
l95Ndnke7D0rzFFEKL53BYXnjICwnG8clobLz/tPFWPRk4qKU1goHkxw7KFigAGOJCkQH5ON8pze
OdVkm0jU3qpItxWWKcYOV3adYUpJjzRTXI0rMUA+9kwvq4OyBTfEHyX7gTyVb+yWHzjmOO8eZmHy
jS/YKB7jtng/uQGErNSQbwhGdqympWRqm3ogA57YmnJI7c1vDt9VUEfQ+ILn8PnCiHeHXdHFu+1s
08CsA+egQ2ZT/cfu3vk+npSFNN6/BVZBQGXX7cEX5jTfSRJYwjWpX/WlcXgIhgsW6IpwrmQdzbSq
Y0i/MIFDi1Q3qRGwbgbvAiryatCSXOPwBS/dkd/0kKMhIVMWU9seQ8+DCCA4cVZdUddBJrY2frDP
GvU/Hti2EVzFCOwGzXeeflJIP9EmSuGJcXgJulYzKQO4a+4nIe4EN5CMQAEG3vXNzowcYLORa5Sq
P7+UDB5gWHej+2RpV8cskRy2Wf8gGQWFXI1Xyas30cKlA2jbRlsAdiWzg1sE3o/bpEqofI201Mcv
kcn+3kLtkUubGUG+zq9tAO4uBFt0NySoWRghknCLqfp0WsoQISIh06GXTSdjspHl2F54BcQAuhN0
750hbMeesN/Nfg0eiFviT7vVdPqRgrHtY+AU7K3tBDWUkDce09/bHxYnmSOyL6WKq79ZdKeBgsTy
RC5CF8feaYJADd1RCiElTaYHP8PUBWQDNYCRBIu+pQHpLrKI4IemJ5HsyndNiF+OEE1QEIbPyfj1
hdfwP/ZlnnTag2d9dQgCI7QSjuFuAVPbHab72JzzOL2S8ueKDGLmusz9ettkxTTnC+CszH89fouv
JFhIaSYvjjsClGdZ+d8dNNIVSYl26T0dIQHaAbP/4+OpquixUa7PDiZ+3YtGnhD9WKO96BcjXwDy
/AkRYQ4+aht7X+mDEV6DcaMvCImnTZ/W8BrfZMS23fYQibM4KW/rfWbdKxLEg7qXNoWk/dsSl7Bj
Pl4Gd3sVtgoUTQWAmbPfWZhkShLWphWdWNbKguDUpFeVw86itVr0doMJGyddgqf1Pj0Glgzm9zTS
ew3GeXYj6bp0GBUBLzgpQIBhKlrQidnW+e9Ir+eTZJxVWSmlCsl8f7gPVPTmXk/2wUVSKb3zguC6
6zGZWEM36jthNIot/HCp+0XUk5IQxYVtV5V7sBLbOEmKhPZOosMBE140PhsnOBKycpDIwVTYQ6Rv
iQYfuHHGLcJYOgfTNWT37GS5BqqNVpOYvXjukLnxvdNxaaItBE+ug42EMgj0x+gIR/dWKPfEtEFm
+qbDV/BA/iSbp+9njKhYUdUdQMfFf5XBFCj1PrWU+uqFTvW0UMEMdaBK2lr5Ym2EKve/580AnmMy
K1A/p39/n6wmcIpUwDTR/Rt/RFzuUmX+2LrSEg7KmD8MKNYmdiSDxfy9e7MJCLsjaJ0rKPqjw5Rn
6rJI1qmy5lE0AxqzFirDAX2TT5XFZTaq5hV0+5HtdmuZ/tekPfc1xR0Lho4JHK+E7q4WzOH4Eni/
76FnulU9Rf1HHNELgEDLL/eweVdjZSMYweo/axU8qKkjcSAfeo1O0vMv1O5V9FIDO0kDIzWA/J71
PGSzRjv1g8XU8o98RkzKM8JPjN+H4JQ22eEz/shO22FTy+EsfVDrmt7mXrpC2PLEc9E64fu6FT6Q
Tc9ADYOo7QNGWE4zJ0wa5KGtibZK2EwQ2hOcVarpcz7+5B9jxkfTzWYlLUAz4NaXL1mVT+hyR58F
YXWEE3EwuCaEydqO1AF6oKcRlf/5jquRZZoIO7S6D0cBs6RiqTEYluXpqvz3Vl/2VNITDmDnwwbj
4uisgoIi7Rspy0VS1qdFwZNDzIt2tYK+qHIWdgid09ofNIeix0CwTZc0q/pdIjC0TlTWMkETdrZo
LOMo4YTAS33EwgXTsQnj0V9RA7guC6TuwhpjxOtFMlA1jgmklxyyIXGDl02pMkXvZ94nF67tNq5E
rT6wW8SbKcNdWn1kYQWrxKJmGFGcPzpeUGgz7kxk8v45yKYCrY9Ydfng3Z2UxAUGR+It3OjcEMO/
k4vS38ADo3QDaFOgxouMehKrFmHIq9nBfdlzFgTItUSRphC6chVF7WOogMMwZEoXmfA7ZHiXL5Qs
WLGfrxEkAzGbR7GJI6YnpA4wgnOKc7vbHqrkrwVGnB0ANYHPLcVP3SQqsacPQXblUOZ0FrBlAxfv
udBT2XT7eNYf0p4xst1l172IY3I6+86CmQHyAivkBpHEbhJ56cHvV6fR3q/eNjIht1H/chsMkAsP
kEhDc5CCZCxBRLJ8e1OmGUiBJiiNIXWzumlfshevzA/O6bxXZkVLy5aZJnamsjbcpapAkuFdWdsZ
oNpMC4i/awn0mLPdA5upM1hUlO2n8Mlesdoeh55ODvmuf7kuk/tphDXpf4oSgWdRxoirIfe+Vew9
3Qy4jJNQJNyxctKZ8r+lcMD0VGk9L1qY3L6pBXwMkL0S5nj2HUuCusyF2wlJpzJ/ST+cVGFigv+F
+PM1c6YF6JgLKIdtIaBw3eTDmqnA/jnfH3ZMs+gcJaUhtrjL3iZm2hZxtJPg1A1Ufo7ZFo2PfB+U
DZU/P2Y9anrYrK/R8KDWf0rczlrcK6vXyfNIkVuPQ8Oqo7ssJYKwvNqO7sB7rlKJnfPAQi4Lc3gb
8REJ0bEosMYm8Rm68XbvnPf6z6AcyReQ/PTV1ulXeJmtbyCLkZPzA4fjg2+Pxyc9pq6nCGlwmePN
gmz6O9ao0ggGe0117ZXX5IxkrkKNE2mPiqWNxnryGa2fs7W2pzwFMlH0wIXbh4xoAjxC7V6swq+f
tlyQ7ty3wsraHHlyq5pf8fZu3Agn81DRHilIEk8w8kulK7SfHs/QFoN7Pi10MOS2g59sHhPRZblf
7vq01MWyjyX3ycTLzK38iTyXTq1VO75pnI5BVg+C3wz2I1z49gV7Bt1MO6VoEnW1Rgs2uTRvDmMF
RaQ9Hr6jg4XyqyzzXpoAcux3E5p7bTt7PEFCk84G6P9FeYWxhS5TITtrf9ZA9ETy9Z8Wk162N3an
UBc72nztSpf6R/WsPQ26Tqm47qlpQUn3+N1seZTwqAKtCQ0w07oxM6RrGjVw0jJhwSB/4uLCIfaE
n+bhFmjKMfj19MNeJzm8Zz6TyRkjlEBx6HmtBAEOgqkzXG9xH1/MIlLKu4iF+twoAmbOyzvA93C2
y45CoRGlos8BCtRI9m9FI6pFfhW5jS6XfQmwMwqfA86/9HgCmdM9M4SH02YxocRyF0OKwVKsdyXe
LIZ7Ml+ZhIe3agm5viRCHimwJWwZR8jvNp34/HDYE2UZGh5Kh6jHk1W0Tn7Cf0TMmZmY8fuA3sHx
4XnpvlBMaN/7bc90mM1zQimEQ5tCVMnNPov1IXB6h2h/j65u1H/l/yHxd64ThGNjmPXEY3PdhrJX
PEw5tT27MPPW8hO2MjnPSFTlXtEBXdnpoTxuNEeThjP9wp6tvcf1SH46ixSKjdoIDdUtmt3onh5U
1UUsVeQLrjDDerHaapmCV4YQuxUbnX+45QTXCrvuMAmTDSUUWrVklbUju6Xuv2kGoQV9djVTl9Yc
abjJuy0mtZKG7hYrDZDqXOA4tYbIZa3d3jwO4ssEa2X+beC0mOtZgrg0f+Vo5ua5hsM60xDLxQ44
2wFAp+OJlh9628qDOSFMO7KyHSAl1dtrXqV1U+KL42bw2BbsVX1DbiBVK5lCfEklrkFHCWoKPuXO
gQ3P9QEZOC8NpVovoPUcZwc6KGjzHWdRc8eqZvCVbLPLZHMPQrkijetGzFTIt2QGKV17mTyvs2Mz
20ajizO7LF+V2mqxZUGBmb10jj8PH3I3PeiOyihH/Xte/JMN17Neogp9dcoEtsB15r2pbyeCHSso
rZxBWHn7cFh99jTZ7snwLEjxrAk8aHjmYKNd8BghG+alp4Ftq7VmiEgvpxihpmW2AQ6Z92bHIS+K
Aq2+QdCFdlkgEhH605RjmYV5AJjbFZEjO/35vA3j/yLLp3pvTMBkfUkBY2HtH12zgZiieTExjHF7
OYYD4NAOLudhvmzLPinXQ7malODU3tRIUkMHBMT8k6BnQB9WXHT5nXtHekB1XCIGWsB5YlqzSl3q
5M4Pp0TE6dfunypboy7AJ8NlziiQ6ZpoTNathJQRn/IO6KkoCc1BbHWCnRbNXNwSIjw/rDOMsX0+
L70GscxmRRnpxGZ/ysbX7WleuZQtm2x75f5e9zmkuDN/WCSS6i+EQXkXBwxiNRI5Lq5PQD4HItOf
N/9OjRIqSwf6F+fz91pCJZQygdOJMr6Ei9Pu6CNcuwbB3x8tgS2oK8B6htmGV+3Vkac5Qss2oESP
ZD2CY4RocGq1OIcjtrpkixxnrpz98hzt3X4WHj52KZMgjzoAlXc93L+rT/4IOHJigX+XpaSArnqJ
CiN8+wg7zF0cTC2yeIKSrhf6rndAaxWCfmLXFbigJ4QiGnx2GyIQsea0u1A2mTkqOphQTEMQmvIl
WEZoNdeke316UEQGLgeYsLUTLm8JAyz3PfS8q8Xu0XbnxPsGfCCbGn2ph9XYCW3rJGLaUlN0zSKf
jQfVUXjj1hGpO+OUL37ZLZa5CrdEIwOH/TwSEXlEpo8e0Wmfr08XMx3Lko7diJtSQ8p/6rbn7FRl
XLCtn6ae1WibYSFcT1WrVh+DayA5f3Psk2gMdH9Y2hlPEl4/MPxoWN5uhLOFE95OkWpCAUXhi4Zt
SJdImu8y9SQCbOlU2GehNUxEtwgZoh/HDVEhOc9dcCVeJAOa672maPMebWB1OQ0Mfn8j2Pr5XP02
NSxncRjprZxzq1o+nCk58fUj2HWR+p9Smgf7W0u91psc5MThk2gbHJFj00jk1yba23n2zz73lPm+
3dufSD2XFVTT8iQ9qTcJrWT+qaaNgxaLo+AX7VwLdukwIY+SsfXXsrQPNIaQlKkY74rWUI0aJSPU
O0RyrNuHE2zoh5TajDaRW6tOacrdtAPTi0tpXS7NUY+RdlCwsOv1navUnx5T4X01lf7NoFGnGQtE
cK315xlvHLCzUtza/z7xECrwkbwtNQqOVehTe7lcoFb25SSltxBpDE5jS9h0xvYhHXu6SZNgzIUy
Qa8/IoWgP76ykQ8ymKcrksibAQ9MZ+Lrjaez7D5xnsLckl1WYUvfIcrxXV+xUwT3MSLr9UwAVB6f
OyM1YUnnYua1YEgKnH2vhd/6wLfUT2VWRA/7YzYpG43aLg+qXAFhtmHi6NXhKXgbOmFwbaEU3Lae
j7hbC7xZYLjU/WBdfRCXTbGVndrTbeioePvBbTBXFVN/gceSiynP4RQQzbGzXjWHckhawBGDprch
ojw494/25XjEP0mEA8rkj8EH7z+usF3u6tb+Xl+qCiUyESkPNJrMVmW57FdxOMbnMzDY/kMHhUy/
kA2fphwyywFG7L8hW4v5HmwRSIkhHZmGW0zJ6SGPfsP0/LM7wcSOLda3zhcEJhEZEd6WK5VGeyJj
20d6gEGS/mR2dFSHgfxQjVOdvoKwBFBKVt2v2DZ/Lp2Mv3KPkx95Sd60PcB681QWmAKc8MfrpcDy
JYbbt/C7fSWvIbdW0E3iiclq+k4ZWfWbW9rCBHRP+O7Vs9P8Wqs0dxqjyPfLpuOzFBZlfGjizqlU
SG/UI2CCJ8pq66lvVft8lNLm6IW3uxpBaEknm88fDWaNW127UDVG53w4LsyuaF4p74ByEXckOXBs
6exNrby34Slssx1YrfV6m8lDLBDibJ8EhELdQLQqheNxZpIfrPv71n+34QIw0w5BLgel//1hJ0Z+
+/fqiAv+wsuBFMkdsSQpMuBq2kT/jTNOPIIREncMuhkLwQnV/4TJqf0rVbfyWoi0UnpF+8Vyf8Wj
9IwMlWLytY8cIyorWy/gwh5l1lGe+AJWupWabqTFQ2BtoALjVe8ckKpmtWvHHGQetUvoOnynWxF7
gQpIWz/q2+3IYRomigaFggyAqQOwMNppPOhRrhrfco7bDKUh+lZATX19GXiUhlclx54dG3XFpK91
THvnq5+IszdBP07vtgh71C8TQiq9kerFpCtQK50yorZe4u3favax+SlCBaRIf1ZiwbRp4Z9TV9G0
E/KTyHZZ5jEUvRWtwLGwM1h1V1Rg8YGQLmuLrYdKvL8yv5TFwfSgBijWJls5VOgv0NeYCi0QIkQl
dWc+JiIyEd98o0tmCxS62oV+IKw/sFZz0sVN4LmrEtBa4Ztor8EZdCABiVO5AdbUGyHq2V+oFQ9n
mJ8o1GmLT8X9r4QLh4Racvv4xxRlumgQO1XzuG2MOHKVDLY+rR8MSSex6skM5v7Q28DS13hw+BCr
oTEBzktfO4vZS+kmUVIkzpup2ZUAzb8FSuFHshrG4g8EYAXd2vlxoVU2e1HSC/5NOG9Frgcx5wy5
RznbcnUhmDUMVYP1QLo56JOyk/Hfsntoouz6tw5kkjv9cUyvNhzha+btIwZxytufivkIQQUvv6tw
o0BLV8nkM+IdlMArsRgmz7TPy+PZ31Q6Qu8jls5zFHcTtewGz3Dcak27gp/qClJ3lbLihJkldjxP
kSDhOLOxMv/yDm8ESjR0La86Ab8cX6svnXfZBUEoFuezBX403vmI0MMEJ/UOFYF/DdlWvn73XBhJ
RrpwHre674+ZX84YOyz6qvv35U6hYTyxKyOHuXVUk/7tHZhOVsaX4drdl+W+vpQJRmaA9gzHkvho
BwwGRS0L/WmmlAyfWVjmPQB/GlmmHChGB3X4FSCtWC6TUk8+chyUQ8PVlb93Z7i/DrDirzd5WFt8
+Jo9JQYVhE2KF46hxtVdMOfaqGcdpFxB0sxkCwPca0fOF3vFr65WwvrXsKi4c6XZgP8xlpms6cxQ
elXfdtdqyY3xBg/2H4+rGWjKQVkQ55eL/1OHsMG4iUzhJM6reWUc6aZ9QgQ5+WTAUxIUPtqqQSy3
hRwaJIuOUvqh/050lFjn/Y4lRRvkJiPuPr/ou/zJQjGNSiEcLX49tWjN4oU/qm1GXIM7n0p9vHIy
Uivhh/uwwyREY429+BKyB5jBP3tZr+Zazc2dxAOrYXVGLoBYZirnbvjVULC/ZF23BrSLddHiS52s
BvYRzxlohPx+z75ZDgLXZ2aBdla/ukrxDiMo+Ur5f0sCXR7YrJVDiEcm1aWE868a9jARMZ7EEqkP
r7pBfT0td1c57pacKaiIUjQduUsbdVYGNGV2jpvXDKDepckbeAWOfOlRp0SPsGzg/3YBu+2TnPCm
/VtsRsrX9PyiL1OpQqAQf5yl9d7duO30XAPFaJked6KxY8wTSgEX3Zk+Q3pPR4ssqWZPorLabkiZ
4BE0cfuajdsOzxIRrMsVHj2W9MpFFiYamlrKA1rqLTuxY0pNor0WYezfTHH6mXnEkhb/BsqgXsK/
FPMJBp5gQR92/24aoAuFyTE/+6R/23VMTU5TZk21M0IEIhkpA+GpTsb7/19PN1y/eJELYd5R8t62
m2dS1BSm/mL0zm55yLM5rdJHAUXf+pXEMttVFis0wTwoHTyFtrKK3n2a0fKiozjz3lTPdu7mAQCN
mTOJ5e6fx+2EJozYObDS7hTilwd/jBjFBDJofj+ioE6zIWqS02dKvnWQb80HjXDmvD6WDwdBhKLq
MsusHEnvoupfr/nSJer+n1EQUqierSihSRI8M0APPXhBAsaNZVaBFhEK/1KTV86iQ7qy9TgkYdFy
yVd+CxTnqJ65O1cHWCabNPg3TsbWcJl87lVZciKBfDW8BKVb4hzD0iEFL5ahjebcAMl1PF2pWFlH
VL6D9aUVnDkiIrNeezqLlHYFcThaPmmAfGbyR1UYpD5HpSDOZ7Mbr0Au+8nh1KdoE0V1DzgyVC9o
RCxz96/37r4nHoKTISqWQRsEvDuqE1HOR0U766qUvHjqWFyFa7kYkNhaarskBJ8KwZg1r5ezajzv
IGGIVQKxW6IuF5TMWqWzOjKfBptX+uxUd0IzZCxY3OdVDHO0fow4qN3jkDJcCf4fS+ZQmu2UmQ0p
XSrhX+gCmwLf0UJLXH1HN1a0CjZlAQbDrpX+BWRnXMNXKOE78I+S1+nS9f1M5oGCU6XV/VUYsuXt
Bv/0VX0NE1v4/KqSHTwGIVqBDwIX/yhQFnWkwkAi8Kiathbbqn1+3jh6e0bdYkGoxe67COgUK4Fy
yroIT9EHW16cs8EAcNR6QKzv7qDQPF1+aZxwc2GF/iDu7ojHm/NabPez+qkHjkLtMOVBTPWg6eT4
wjY3eXYvfNYx+K2cFAAF2wN30ctAckNK5teO9K9VMgZCnf+rjtQHBahFFFY0yCrhOwsqtfK/Mrlk
EykDi9xhIUc2rKdJzHPE06/FGujP/bb42yle+Wve64gzr66JUSac1WUePoyGGh8Sak/IMwkgKOso
ySkhBEdHJS3ZNO9rQjDFOa+sHmarxJXH2zhxGaMqdHSe1pyHO8UklUbEB/fnrTHqy2pdikc89xwF
U7NPnFTtTO7vb4FTAv3Q7Y+yDQAev4uJbsOdfqfebQRa5y5OmYj2/H+wk/I3shxvOQvM68FLSvKI
7nU/JH0BN+bkKPsQYV4A3Nq5SEZvYbmI6mlEP1Flzov3f48iRPyAsb5BBH+PxNaAiN/hBBuvgAmF
vSVgF3aAIBZJdKh2FhXJfYo7/eGgZ4dwIYSKZ26K9OqZExtjeBcc2mZSWt8Js+13rx6VmzeUqreh
cJcf7WIBg9RisjgTG39GCYRMaKJMciNWQD7g7Ik+eJeQtiMI3VtqYRKLeXQ15TgTAwIc7OmeJ44p
Lk6kGmcw1jl5y8PkLhJdeFUauvPFxTIBzbcPMxSBQmM/3GjmAWFx+Uhl8ukB4mHphpTd/10C9Uh3
E6IaGav448yDOySaTPtlYOBi4oeyBp93gQuNaVMq10bSqrzvlTlxSo0aYj93OUo/3TwpkWJb/lwm
m2SfjMJQRbCfOt1CifIu0tnHjPAkHv1fuYlUQpajm0lx/QwcEinKp79VGVkFHpA82ItAP8VYEwW4
slSZFo3rVM3ZjBHbHl0E9y5EV6LdbBcdz68/WDl6ZojQdYRAAD7pnW+kh/CV/GWwgDyoR9ovEaKl
ANqmsdkgDKKdBsmI3VvERHq78QhJrZWTBxQhNHo93j0qhOJ/nZpZvu77e/YQl2sUfZ8AMYKhELB2
o4arMVP/gcAm+pOZB0Fp9TZWXpOdG1utzxZ5Cc5C0jgZywgbCPIujB5/d3vUY6WEo5PBIJJ6gf4G
KyhKK7Xx6xnupicVEVz7GeOpweAhVC8nf3+K7fGaReRy+/idYIThmDpMf+MhcfxKlgf4sc3WDwSG
X7VPn/hnCAcA9oDEDW2gokNKQgWf9g1wQr0OJpeabbFaRxzFmukKsqEt35U2DaIEb49ECyKRXndd
mXV28QWvok3edyEd1MQhoHDKZns+QeT34BOH20Ug5iDiMNx6yUQj/OBmCt+tc0yrK2pm0723A75x
+stv+I0aOA0MwJQLvQBfusGySvP4gul6MCRDz8p90CKmS26ThJ1yzXHhOth6l21PS0ifakNVJVZu
q8jRXIVUYCnIQJpOJrUQiBY76AEZu417TfHiboVezvYCkQ7Ky8+b3dhnA3bLqkgEvOgijaW7RDDf
7IWLCQ6YdWIjWGjzr4o3LQ3WhfrY/IzRRCgaQ94Gq5f8kDwHABfD9RqvtBGduo7ly04JDXt8FsYN
j0VLyYj/hdLTB+oA24dP6eIvW34UQ2uu3P6MxIA3zbJvQoNYCkTtgWjOWUb4k/Y1bmygWiSVzDrg
rT8ZvCQefCYMEh7WDri979p0YGu3ONzTF0MJD35kquu3S0zylZX82na9Qhsm/Gu1CHqjzeBpYeyL
DrqSU9q3mhjHtDu7OCNt2TBEl5VKSXtUS2XEnQEBqdhfSTmNBQNWy4RfbZg+qTLNpooVzQKhpwtI
2QZx75srr3hUX+7mq8+BRkWm5aUjadGoLHVCCoYc1Ds90HQzLTHY5U2elnoUBTf4Xq7ihqqPjL08
T/BAKPslx/CtBBkKMr4RAvrcj/RM65icv+tzrLkjBNXbs6nppkN1IBkUEL5NBTwBGsg0skd/CaR0
6p179Lpuc4Y7K8i2HjyanOKYHgV7omtyZXLTGBcEkcp8HN4kzHAA0z2rz/iV89zCxvI5QQcY8bn+
WSWCXU+U/5kfUniyIjYDqx0CmGAbuQVSHLQsUAxTaGBmHR6NzJltQAoVlzCldBiF4DLmNX71LbjT
suIAVMrCXLr23xFaPJzCBzGqthb7m0n7xDKBy5Olm1Vn/FAV0UpO+2QK2UD1l04yvEbIrFnGzz1/
KbC1XrHuvLESj168ehvdEcr7N0/HOaFiVcl/Gj4uqZ6NR0bWJFt+m8ysG1TemaV7hqEuW3v27GLe
rNe5rOcquzn1NXMJwtYZjswxSdZRSwpvA9oi0ppImud33HyJG+8aT0AJS7H12rYUZW69vDtRHUhK
Y4IitG6AFOCn1UyDZmx7dWBHA9OYJOf2PAwvB/KN7aLZYKCkazEnb8s0GYR2WgbLcq6zgoUegPHC
ygzBNiSH5rt4UNQkp4Gv36ZgnZ9nSDeYkjVj9AHg/tL8Rpwga6esdO78tFC/I+imPFc4Ow1BKPUd
Kxkw6n15T9dzrzXFXD/NxtkYzodyiauyxnirsVlDqbD/EnS6rbSATW+X7td8RSZgsLaY2oGN1E4g
Pcia0/umFqdYF8NdR2dv4kDhH4LBfSMMZiNGvVX4WPBrmjJ2OhJudtb93HyyZw4cpXJAJZhgJZRd
b77jlqo3mXE2WwJl7d9tJd1ORKYawEfwPLDj8JU5oiA7wpBwKROkQ/HThcpfKvPBr+ZdpTEG8raP
+GzBfwiU0xjMsisaXl2dLqdvO/ZZghV4/Z5x70HLP4nTyr0skzuLQwPmOT+lvVVD8L8VT31eFr6B
M2Uk7XlNNQn4UXsV8tgCLXJQOGJvWXq2ReJGy43IkVLuyi84K0kql6/9IAnsK181icJXlP+4NWNl
SoQcDMSV4bWZ4/VnHvQZMCHerwV5pYeRXMTeeXuNvr5PXvn/Qvs5gYHjaxv15hSXvq8F1P+iqFMd
xi+7bwSkJgVDSkWJw8YBhqIlHknCCneE9qUFomQZNkk6bdEc+8nsWVYM7EkoD5C5fyXBlmlJwJwD
PGJUoTmjNQZXl8QGyqoEBmiACPP92w4VIavPsKfT5QvGgyGNK0Gs22RenwmeMazHKdXRF5rQUPGf
Dyh3Gl0kEUGFVV0WCtSiK0nHnMorWmn8mF3cbUpPBB5HrPE8GBfx9pIMzwN3RsUMEY/4z6qXhiEy
GLsD6bFFFbbAC9guTc61I/AsgG1fXtN1XXTStZrNA97SQOmhPJGwQ5Z1fdFPI/hA3WRT8Z3ssMmX
XlGpZNmMZkdHofQpEZp40Dfg9N6wnWIPBOjNW8LBAMYBNR3Xj5DjINpxo23QafI48Ekfi3BgKIYq
QVWw3KnYhDoog3FoU65U9glN+KTDnvSYZlO+siDjoCCd/YYWeMXDQMxoMqQp6ICKk3b5S+fDs/nO
ziKVqGMQCe2S/hzjnfsdWpOaF8T3y9fDG7ycvxRAfyzRAByMgSS4OW15xWO3JGF75Pdm8tD+bkH3
nDUf3z4gdcc3TEOby1+0IdXOXYkNyPuYSaT+qiYqvPPq5HeVZCatJoPOPs+PrtvK5z5ln/bdj1us
uQKYxXzw7xxnoIiMUUSTIbME3zGLyYCBpx7/8I08i3h0PcaHyZbpxSgjNA3WYCuJJMpMCbTw/QLm
81En+FLMB2Kn0hdYvjOtleRgCOzHr374Dh1oP/GqoGSd4g8TZMHnFFNXensbE4BBBBcXB5WP+pXO
jIDrEkcLSZK/q07zxgyBNoF/9Qq+24aJ1mSYUUZMD/C8ZjmEqC26JnFI0ymU6ZNgelSEexIyFc6B
cE2XiqKv1SdVliL61xqD3j6yhvLpA1O+SwXU0I077FFeOAqGKPaWukhfOSWxH89fUxQbi0tHDNQf
BHqkmDdjv162L7ZesCV9DMi/q8r+zPqVqFq0EkG8Fg/AGKy9SLf5CVlqOg6yXeJ1pB91TzHTvlYN
G6bcsaK2Zmn5ibEkRbD6EVeD48UHca0rN4D9HXIsCmX4LkstvPfnun8mPBTcMpnvYNp9vxKhVkcd
cHJp+1PRXLtIEY1wtZbHnXUU1OEnil9xJo/4jR1mEP4+oAzzOLgSKtI70zL5K0W0e55yEgmLDjZx
+UxoLu/NkKeENnzjlWeqK6G4Alw1hiiCObbb7I/kV9Hp9ML90CLRLI0gfvKF4YoPBTAsCpmdsUDI
ldoCEaG/scgCSwx1d0YbbVQULwdqs+e+rFdJj/rxF05meFHVAv5Ao03c1ef9ogPt0MNqgvcGZYCp
7Dpgkei6vigbcnkIqfgzzJeULzzEBauDudo2DyZMkm0VeoN13MNLiUhrI5piUp4CMow2YQFlFcWE
nGvX6NYU0+CS1NKfOu5iqntoQqAuVNdRC/NtGVR79tPJYvkBF7dCu3i6fRK9eO50ojPlLJMyW1xm
f14HYl3ToK+MaFpJzJqgM9jjtN5uckaJtcJBSA995W29DNcbJffwOUxV9EfcpYQqkN6M2X8DlyqJ
Vi3jS6kparbXSlExAbbj19n6UiOj9PFYs9lC+V9iNUFQ3+mww+jAhWEVmx63osE0JrvZFDmMbXJ9
s942BEwIYyq5p8LChlCYBjXV+TeTArhJjRsc7N5lpcG1yRlksCpbmGRe10AgAkZEw3u4VsLWqePu
jXOzhrs+xEHzUWz4NXRMQacs2tWeSxMaEhRpfGWQR35tk1y7NR5Miuruql1EvY956VlQT1rxDXMm
UpxmpU8WrvC+XOmbVfTC5lZ9dDAS7gSAXvVSSvcjCrD/GbdUn2iJqNxb3aPXDjIss88VdlGmzfVn
9HrwUFSw3s/AYRhgdsOIBOMzyR8Hw7FW5Hn2y+wxaqeozhPzsGVNij0izFLkk89KxgI7R6HirsLO
BFAtV3pdISzpLONqZR73mP8J8uuduQ613ru2rnLK3tLU7i4k8e0KsNJaenQU6P8jborpxfdCuUFc
LmhMRoNqsKFSkUunR57UkT/D2fb/M8Y7MYi0ghJPNM1I6lDRO8kQ4XbOBs+K+Q4caVfu5L/2hHT7
qJK4reakOYQxKcp0ZdqZM1CwVNrxMLcfn8adBZIBlwrdk2MNfWSc8RIvz7/g3S3JsR+3tr4GWloo
JugaklD6fNYH9NatPDMqSfNCst38ZsQwdMmounV6NWJXTDgywZ1+5soCX93UO/kgTozL8Twm7QaY
OpjI90DaL2Ki94a226vP7JIT57RSByykT5JQtF5TfoLT9b0s7aHEaCgiDfw+VpIymHtEBxO/kspR
VnMw3CjwiyrFylPKp6gk9J6sNifzBouRrHOid9HYQm8FjpjqmNV8twWY3NS9CjEDcqwwnLe1uQdW
gvshITBIWw5zawPxqX95FjrL2hVFw+S0T4by14b2spQMbq5v/GsmS17o3wSM0WOLY3U7+08FidZV
5J+ceYFO5Bt4ZEN06KJaYYP0I+Stpo07OGQqyg2QSjmttoTWz6vD4YrXHAmfPMZOr4APSHxjKce+
YiG5Av50YSdXp6b/CuEsu/J3f6ym8ndVct+yRzeS2AMyR0TIJZyLPphhOZowK8Ap52ef1arWh4xK
WQUjJTTcdPYyDP5qR20lswTI661AWEgaXAwERmVkq9JgHbOJSIeQEyCEGx/JOfv+9GpiwRqMiQ0R
wWmN7qib4hTyclAWZCTWytgA1xF7ZRSiyLRXQEgEtskJ9QMrV5yS5UdjcE85OyoT+s96okRT/AVv
9fPX+6C6mFo1aZFcE6svww9QWHqaxxiDNB1r8bPjJm5cF2+oSHBmp4G6dl2YnBCe1Hq2hSg4pr3s
KOe0vGNKmcBv1XtjEpvuL9uOx8rdzI/DuYVQCRSNplY/bVRfRMOuu+t2z7dC6Jty2s0A/RtvA/ra
fDDDFnw9cfkK7P7ZVqK9vyatYwvj+X6zsHylIYdPj1E7nJCsCTsO7TX/DU1E7bh4yW0YPakkcu1E
WMsQxu+maQBE/HL5NUCc42Ee7jIE+sFiYMat/YR51pK2XGUIIwLqcXTOnKLStZ56KdYs7Hrzx0IK
Jljtq+9wOMmuyt+afbiwNiHcr8YZgp4eLkkaeg99mBkEzFu20oRK32JD+tFXrgcehP/D14PpZ56V
ueEnwPFeJ+ROk8llkzFf+TX+6mVJCy+csjjL6LFMGeFHRIWKAbBsO/l/RnZn/ObhMN5/uYq/22YE
2ma7/P5XvEYsoj7vQ9lNmYmmtkhQRFOj0Uw1xG7PLH8Uh8b0ACGF7WYAvXdzcLJGt2tB3Nm4j0e1
f66fpsjUcxS7+BCTsqUJAITKOip7JOT2NS4AfOqXD++OyEIeChl7boUgRSyl36AnGYECxgjgCMsD
Om/c+WGKbZEjY4I2GpIRB4HKewIYPSRIDGqXwtLlz19TL6AykDTaLk6d/GhmMbKlM2Lu23ildRQU
vxCmcI1s3mg3KZtRUmkMZgMDpu/ZBDLwPGr3Gg9lzyCAR2kyjk1TgfKeuU9AhrdXoXulvE8rAnEY
qjPq/9hKvOXw/Q8Yd8ehEnKMTbUnFSC/15aq3lFd+CIqVdxWCHG/P0UhUpErYmj73uL0CtLSgmIW
73tImR0XT7gKVlSKo3jh8SQpzSqkpuOj6qkG7QJgr8Ch0OiZHyBBDmPJu4dx0EqT1XRXetkZz2mM
HirwjB3cbV25FrLhbStsSwsqDrjHjvbI9arbrq09Uj3MaLyw4aPwbIMOzYBhoBiJ76WHLQOHogAt
jTIYgJOYimNZ84UZsI5VxUYpvNl0bmo1Qe4o1frUXLAHi11U2pFN8k8A/wM1gLsQfh2i2C4Ewd5d
3lxLp5Ogg3huPTSHrIEMSFFOYiKuezv+1V/MwO3H3fjZy/S45nCKKTqwTY0FUo04k/CehR1x214r
HHaJzxvsRWV2IbWvm/ThQmQ6T+M9c1/v6wes34xReboMi3B65seLV89H5Ia9fW0vWBzAJZLvBT6n
P4Kfj6ZfnGVeveC4Nf/ICkZmo9JU7004C3dNhyyFurL+tt5ZKafvP3aE1KJ2hCj5QvZNdpkYHWAj
YBDlDltpYyhbaQfaa4OXK+8fl73wOgA7pCwbu3na9vqMHBhZE+xTPO/OgsKwqirZCflc7V2gJa5b
kIgZn6bepfEUzFYL00lARCqKIk1ErQCK6Q6FJ6xam4Y057KpV9zzDv+/rGBTCTeWaBrKlLblmkKL
jNO2/j4AE3LR3DyRPOj6NBVdFWCP+Tq0EN6BMi7zgDDufhvEA00Gfd9XcOuMZWOCVdnqpy1ENjOt
huP1M+EbLHr6ngAH+te1brU+Ekoi9Br92czoTIh0Goxnkz5FT49r/wEMX6DQMQJWot/WtxtHVeP1
3BcBmm/2taJ3nW9DNNf0YBMI3slIN06Y3n1doVJR6maJobuNTmHMIeInbQN3GKC7Cr48EMrgNYij
PBNzw/LeRZqD+sf9g3nhRHDHQLvsw4rWFYikbf06ZbgHN5hVDfwH0z7n0riU35tsssaGDfSxueQc
+L5KhioW8M5wqvUoRmANgKoLll818YEpHN6nlbXhiQjTL1b6PR/teoZoRcVX1La36iE1kHCI588I
0rgMNGz/y7lc/O70wYt69GSzEgQ0GtOgZ+K3J3PkQB4TRR2p3COCJc1HYHLfTvHn8xU0Ii1iLZ6i
0t6GiFu9uD4zthVuc6tkNcLQKQBg7gdlt8xTsNCath/XSEChk1JjJoXC5D0BkT83tUouSH45Larw
PrMEL8EvKy/5PoarhT8TL7QImuYgZTCd5QhoPf95lhVS3CGbR4N1m8PZrzuT6GpwmtGcrobh0rOL
d5yUmoSopf9jvt6VqNPWl9VsMSKl+0ilgaWZUZ4G/trSzPOiHQuKtusk373/JQT8yOMctQynDyZ6
ejRXrowGdvNksBBpPdqmKOQThGkl2wEc/VcLJSQnx7nAENgrSfDP0QHrKPb152h76wlx8ubFB4zD
RUaFe9iPODlHxKvbpw9p3TdnosQoOkI+TSMuKt4kdcQjrwhFU6UFBKCyf4WbjWtGmlb+uMAIzgOd
Sn+Z1XcU4JSpofvd+PMVEqu6a39ae3J+hxyssAazoWq3ZUpovWNXUGVCxrjfEu+HJDCacE1EjRN6
8eT8LRyVtsKCu1DpHEBMqdMwCkfAvP8nM/WrAeGTFHKI6T1mSp/pDDDQCzvwJrHeMPnXwtb9Nn12
XnKTOngkErSZnfZgIW/0qOWvjqdqO+EKWlzNV5sYIStldPtvkpl1zTg7+qtTMwBI67vWg3qMqB2C
INUTLdLry9/PyxMiXV/l/gopU7TLB2A1PnHZzacxiDOYoDQXli9F9i5FxCtbUlLGf/TLj7dMV38p
mDL/BfuASFNDmkVIxYqATm2UAN+UF+3Py9KInxiwCFv2ZwkSyhe+S/R4dJbHFgrdAV7+ygpdgZ6O
hxCM5Idgb5rMLxlVi7f7zTuTLe6KfzYF0pGiBAnwQ2ppsWkFaqg784vAb011iGMd0BMvLSahfPBx
wa8Tgno3O2fMv/v7kOIpCmFNwKhy9wBD2TIYebFGV8j//q8EoFk8s+j4j4y8AnemN/Loids2mhvd
yZa1/H9K5/U/vc7uHW1XPFAEWMfTUbgxi5aWn70dMK/mkFFpXyqoJVBfdNKH+r8tkPp8rFeOfQFU
izkpONriC6tZ1wlnfYNjV80jrCEKXiJkX/Op4oK66+jvpsYCSZnYyy/4CohxU/YYx0hbYH0LRgda
Z8ubRy9fiyP96a4mR7Y9+LPcYZ4vXgNipulIJXM/CP6dNKxMBPPP/5XdPNMwSxaOQzdnmtZuPYmQ
Wtjqp2iMi0Dx2nw3tklApvJ/MQ30WuHNab7VV03vwcMtfeWOZ8z/cFhEbycG/DE/8bVPYhiq5DoJ
J0fhV8WpGyEB7kSpF3e8AYb3BsqVo7xB4GElmPpvKXcxuCoMELS5SizPJLklKPxqij7Hc4Xp73IA
Pxalazut58YSoAOqeslFv8TuywOQFf9a9L1I1NisFssFcUBeKjd3rQRxhbL3uf3fBsV910J7LDv9
LhvHgINhwLWdeBXABpVoZfx9eR5heVCiEcZYcnW0dSiKD18aY6czUz5w7CWIglv7Gr7DuEhCrQYq
NluLOLxoX9DjzQ1+yjBIi9keTbgDFFHNg2F10xRxBrasltfNzmsqETp4UPZ2ftq4RvqnQQcoxCjn
g+AWAgXv20tWaQl/ze4l5NXbEZ9Vu1fVL+uaJWLEdg7iDz542yCCkZKo/Mn9yPrJIigC7vzjFE5n
5ZfuZFunlXWlgy5yzdCIoopssNJxA1/V3Ffn4rJ/m3xoOX1J4bBAdpOGIcB7MNefBzj0374RJUtB
PqxUntyoHYNXkHxuv6SoJFn+b+lZEXBFZIKDz2BEUQLcffMPLUnqK6QEErH1woJ0IXdRbBllxKPN
QypnsjXHdlYznVDj/tfV1AYtinSzGgf490UJ8d+4V68hKmGN+kseqa1H3aoYtV8uUnTqIakYM7bV
2YIYtFWHBbCZHb4/RxbA0nSs4785hU5DHdUlZ4m1tx+vR1pLZtKg8cyZcQBkdr07B1cC15gfJ9Nz
uk5LAkW3UDsyboiArLO/vsozKv1lt3/ncatutqW66cGh8p9ASdjD07ouWSL2YlZ4k5TzZG4nfbkb
vnNYQ8/M7zHi92MQm4L7yNSGDo7Uut5jgR2vBePLUE/OMOGKTuHjIfMcQgYrAgLIefWjNu+bI8cT
grC2FPIu2mGjorbFs18YjR+L7NSQY8dyNyNnqDCrK04I5QFByUpPjl6WxZLVBG6QGPkC9Ukk+Zsc
yYi+PPmGgcHqH4mFQ1UM7a5ZgzPf0uvYgy1DSVsghJDykqi9UVtiMYZF36Q4FZt5ZGBYumm+pF1u
PWvjUthuW9DBAILenDeHN9W+E3349U/29suDpjvNUcdtwAaKPVNSApNJjjoq/xvO3r14thfWGLU6
NjAZmOOhTKpooZbTMmp7EhtKNN7WTApYR0GqsNRShiGDJPB3ctiyzcejnPlwcTUJMnNdo4LfTCnk
0Q0En7bVMBb9oCAthvcl20wXD8FfKEZ46V/DhDf/nC8nfndyrBVkoo311qlpmL6PBZUSiXe4K+Cg
BOuSLeoytk4XJWaSvu86/wgfqDae40VnTK5tiTUhQ4FyMPATW259g12Ludn6FO1yG1lASLX89zgo
KZrf34m67fiITFvUAieWWAUv7/9F3ObRbU8FBar/pUsrSOLHAycNtP8Teb03KdnRK4TkdLz6joHV
hBYgKl/e/pzXOyLbFcCbXaHvNlbQVbFf9ug2wSW1la7Q/IxlbDxvgd3J7Iu90VGnOCfdDcXv0kig
L1kYZQTk3XlcysHvmGm2WELyVgIwcUUFsu5YMYtyUtzEHkv0P+lBEoCgq0jPF7GGQxWixRJQJjWr
SvXohDpyySXt26mwWoLyXBN37KmmRfkYwRzLkB4jh022UIEiibdLaYe9cIcDVbNEK18XmMMKGaqj
BQBDTgIj6OTzkOwR0G+ygiz4WlTtn99Pju2TSR3Qb+PW1wgARUktfV+dzBkjy6IXzqZUskBaL/eP
KbSeQPcKKzSKEKqBF4fujP3/Eu+f/SThL0RtuTrpacIvg9yakFQH7FnJjT3x1iwrk7dRHHQP1hTn
NpFFfvr0R43K3xnzG5N+GkmOmVUbfi0R9Y+mW+Kz36GVdg5rj9gR0VpEz0GzJ7vkP176OSnPDHjq
R3g7h3FJfmKFmkbRJFwIYJAikP/ZjkZbJRAtBUUceX+f33WRf9ynHR6PaMH4AKArE7di/9aUIyRu
HuHHBTdMpZqC89JY1gXBq1zL3lRs3rbpue+LH2vM/MNalhllW7y6iSaVTpC1d0/LXrzhfLJzNf+4
LlVNMbEn3UPGKMXM707vxCRdhoSJlFj1WLZMwrKH7BXJf+NqLaEr3judKDlJOedXD3YWFDNonKjB
L/uOeTHqZ53H01KHPTZJaFu+r5ILYmg2sQaz2ROUHMIP+50KVsUJ5vyO2BKaENPqXzb1ZGfil7lW
i33KFUGKSDyASeaV+YtMaymZJkyt8ciqa6q57fpedcuy7Vhuk9ieseUC8+56ZWoH96I5/YrXgEWi
dG0mXO1D+9djmSBs+GHq8WJyd6hSg29kVmP+4SE1mFXm111zOBuEt3nVEdDqoMpp1IyQ+A/nb7nd
HoRPiblOs/mdrKsYo21Ef269hda/m2U0WMp+wwCnDqqQ35Y8tPpU+TTdq9ATPmiPpGQLbgP/AXVj
p5Ph3fVVsn37CRbW6btWY7yhipoB3IbRh6rGmSQODX8kC6/wltWg7L3V0lZ24KDc7vQxsXvawalW
gjW4+/KmxbULh4UVSiol2dUSBQixtexHCD2bueblOr89uE3NxgkZMeUfcNHuZDiVfY7nHDs7DGUV
AO2rpZ93i4RT0mIuar9txcVFvHomoLfkCvb9LFPcTrAtM2ann61+P+y/NPzP5kZoDFn2BGYu3fXg
ilumrU4Kshz0nVZ7FAnV5ObPav+zFkaZ25T4E7ApUX+SYhtTQtQdoQgCBsztNB3gk/y7DWinv2Qv
EQffjX280BgEySIqInky80wanBtaL+Udo4uaoWg8WXg1IlrXJd9KURp3plCDc/HNL7Rh3LAf/T8w
jsjn98arm3L5R6MMDyrWVMe+x/E8L8zYUGUsz2uHg5jviXWy7ipL3pLDSXE62yFb/mN6fD7ZShh0
fruNMIgQpFvurJY1kyQhDRXyvHrwS8W6dN3pU92TUBUg6ab07sDw+MdlkCYPvnJK+X5F1chUXGfO
f+y/SnboPlMA4Fkz2ylbn9fdAqD5PXcGuw5fjqvgpGBLlTRLYMp0G/NKcORw46VgxXsgdr/eLd4u
6v9AKZACykWQT2wUdZoXgR5CmKLtds8h039OshCd6b96JQRoKAsfFu5S93SDpvRmFqqMTshI4MZb
GqZicUAWHfgC9t7YRqupKu6q/Fe+8q5wQDp+hV5DQTVWjICUMDsz8hHm7JZpsh1un2KJXcauJ/PZ
R5xPlx27kgmsBXY/M3MerhpFXJeCzZB84A7QWaf0Usa+OCXG06ByZEZ26JjkzHGP1aaa7wqLINix
ne1bT4xUQ4J8UPz5hPSFBGHrPjTT/pqvUfBOTzBv7OUgztaCrYs1Nbr74BJyWaAGQh1jqnpdya6q
p+tKK6vd0mUYEH0FOegWTFi9oCta9YJumBrzESNFh3DQxvAzr6bzCwxu3/5DhLf3Y1n0Tcxt4LW+
DbFEO6v1zpsoP/nOYhsyW/c3QB1rUe/U6OOliKIi7KJlZDzA/WYCrATgMduGMIu5m3nmR4r7SAGF
AaqLiXPl1RGPw0DRyXprvif7ypXntU/U5V6Q/9WTKhCiIOJ5ALf6u5+U4JktMgpd/nNNJvaalCJS
PQtJn0b/BZmJYKESUA/HK70acWW8W8Rq8X0lKJJY/spLtZj0n1ymhtOVOKLJK/6P0td5ZDGmtJGi
hgWGIJ8B5mPqq6vJqvPtVhCu8wHpZsvKqs0b76terehegxs6a1ReUxtnZxfm4cvqAiL0DU7LffeM
pPuNJPVG+g6LMnsR4ChU/loOB/MHYkiKcAQO0nRvh/8E2zXgLXQS5Nkuzjoom6dOmZi+ZTOxTpwr
1Zup3utwAVJ3ZarxAnUg/3HvuiQqsLtxtyuhMRjrFrZfkoHdAzYZWoXvMIR+NkgpB6y526Sls1TO
BwPH5gwIdHXNR/2BJ7atnB+GMI8Qt4Ipb2Va2M/h1aAfiyTq6mzKKBH+7k3pn+u2+YKVauIcb11a
5Udr6Azi8r6L2QzPXNb3ZhpeMouPTnYqaK4dSaRd+lgXTt+S+ysW65QHYAz5Hg1FpJTqdvw07OKu
2ls/N03xn2n5313cOP93z3shyT9Vkq6z30GZzX+KIuAmjM8gVK1WT2MQ/abwBFk16tlW/J8EaZw9
Vo2LDhgfKzG0o1eV++OclKGqa2nmfiFu2w5zwumJhEhgbWp81BIcDzwSYRCVNNEs14FRx5x1OQkR
6GvPY7nIovhrg3AYwW9KVJCir3gyvPuCNxhJ3XvtElQYhS5mz79PDq2Ywv+KGaXR+XiHbvKVvJxb
Fw+4GH3OkbdUOu8olpjIArdN/aph5YuBpTro4H/iDwOKqcUNygCfh84jUf9RHQb5iUHKLaH6mINa
NlOq+sqMJL1Iz+ayZLasyLEuddQBoAwl67bA00PArlXNHt8NJXRlRBD1peuO93TffCavHOqiXuat
pyuhL0/eFq2koP10UHeRvJt8FsMf5A+apxskD8UirMMThj+0sLdx9yFuRmzInIO5NWvkAP6N+nx1
XRazFPVnb21yagF1HDn6ITaH3Nw5ePsALRo559zLcNv6tulP635mKQ4I/fBETNZCLpkfx5ZQtKR7
DyXjFuUa13di2gD8u+4WL2kh/tlguKxFteuRl5+WhlCtUadTamGleKZV+VLfT0yB+45gGJD2wj56
G04MzuDO5aOKXT1I6hcZJD82b3p+mOsHkd429V4WZsOCdQC+aeOr0vGOVG/WDT52g7BTBtu4GUr1
ZfGZYzgJrWyHhBse+373cGlRQ4eifh4he6pa6LNTEbtHp0w9C9xw+xxexOTzN3byACMfOO3o+Bmd
CgnE+mXtc0N9tkmGaCyIPB3K7S6X+cd580msqewvt8HqbiO58IN1xgm17MlXBX1rsKzIk8VqMN55
lVLQmIM1IL2RPgdU/0MKLN7hk7c59HSiRFp/CKc+F5rHRzkUhPJGiyOTPFsBlCwd/5LJxt7F4cDD
u1gyRiThDGBOb2g4ewA9ixNYYMlSZVnjy+O6s/nwLOiZlsFEijMSpoxhZxOvoc1mk6Qvk0PpiFYh
WkO52Ds9vRBaRtVZzpoWh/vXtUDgQNRn35il1dpGCKTn6HjRMOJGWt6dXC2GyGc6f5usMoRRbcGg
Lpy+Ii9hNmWYvdpA5jakWgM+Tnwvn+UI52Xt+GkjmCP30zpQKAxj1byWXNhuZZt/EjqGFs0W9keY
BiFgjbAM17cEFwZ66bGmVclpLJIXkLfLOUMn08cSTHDOxeAmxIyBMlxtxzxXzqNqfe2o6pmiv3Ge
aygXWtM19KKWmde5PhIsZCckieIhNoLO8MU5+Zrg+LdL/rjymx8ge/HjQkgl9pmrXt7v+1mF7q+H
ymDabUI3p8fyIF2C6c9WCmB3yT0PR448OUIl9up4YUFLu/Snb8c1GmDFivVel9tUDngDgcmxKJBs
KxPQ53oRZaDbBigNzTGrwG9cNutU51FyibMwu8GqHNA4Cw2iWNDqBlqrk+q85KE//mZd5fPnrCef
B9q6X4cH/SOEqP35cuIEC0fLsy0vX3MKuiLcx7rMK4hjrU8XXQT2WCJdnni6RK8EjcHHncjcRW1g
nvz8yr0bO/QMWi6hNxMov3BlSsPuFoFxCB0k77CwCYMGWEpcRfH5X0bqL7b+bKvbiBtQFEIFlBIA
lz5RZjKNOfpwB1m8ylUJKmSI9JffA7witupAr5RzsXS5m2HQFuSB4OB4MqDt1rSE3vzuJYJbbBH/
mE4TrhF8NOR43Wdm9bzPEBaOlVqBsCHu0VaB2vrOqsbOxnpGlxtsIb++4W7wjFcLhKkJF2021Zrx
KCm4RMrQwQsCA2mPzI+gzm1Rkvo5Vpr+c59Qc63XwkpXXmO3w4zfArWq0/+BV0i/m+xu8g2rA0vF
o8HIL5Y92r07ZRwZD6hoeNO2C9BccjeH0ukme+//nMHVT7cm2SzOF+jrhnkOcH+Rm3wCFK6uQp/a
vIJYS8so9uPqkKdiNLWasUnD5Iv4mrB7NBdYwgN7vHu845MPED4ItJH3u4hcGCkb214L8UyMguXs
ocvxLe8+iaE8+ktqG/Mg4+GE75ROPlPzEkq+v93XTYizIGtxVBnUsjADb7R+HLmRENBcZAlYThNq
RTAASRNsuH1RetcU5rbj1knk0aggF8JrXaUIu80j3GCGfpenB8kxNSzohPuotw3HpoQIhu1HwgXV
HXwBGc8PP2d6aMBRvphSYute3H46/SvwusViuEspisCBfittHv4/sYjOcNuvrLlu83ZisMR8DxLx
VmgoiNn/61hYdqkN/7d1cMwxcyX4qrMgBk75WxDXUuoePVFw9owbSEejPsfF02j/njleoa23oSFh
F7SSlYZqfPqGTPz2IlDzYonZhoC+TzOQXqUzwHasx5mhbJHdxkwogDyOTsOlKJh87lfYVh+1M8df
QeISutwrE8IQD0u4kb2FK8i47i0GpAyGEN+pdw4oI0PD+Z0FJQCWjkxA3MjAtmOODWTiW6ifhb3n
/RyR/s6bUHAeuq1j2pEYg2kcHWjEEdcrPQNf/tdMYYG0KyOwFjt9LO4lGyQZbRi6Ig+uJ/F6/cVg
2iFqrfjRZrojkESxbfjvHlWhxlrKA4iKCyOWu6tzfFigJ+7UWvOAy48M55MvMKa7DOzQAbsbCE7C
xGJpJ3xQw4fcdNbyPNtQHJIYQOoj64LMaUNvthBDjXlFyXJB3Wzdrwk9860ZHMTR+fS5634IrWCh
LETQHNy89esL7Lk4Py2tZqy3fFmVqW4f3Ff/qcM1+Wu6pPbl7Dof6WCNkoYt9Jr+v0Nk6YX0q6Dq
K8dZMIJlUBCMhUU5qV6NrcC/O7GJojDutRteIrxRW6+9lLFYVjFADQZNF4zZmWpSOD4yo0ruA8vO
wGR41LLU2+zY7BS3sRi+sA3B6HP1ABgkf6/5XRh17c+kgPb7eSYe/j+iU+srRfniC+6OaGUqXS6a
mtmlGneTwh5QhYT6NC0Nkn6UjVGrHBR+4iCHeYMjYcJHy+Hs8Ex1JC5k/uvOKjzOPQyUiPZOCWhz
AWjhavWvEM5Gflq4ecPmxms3z4z253iYoJHE+Mbh8ddy66DM+ltwEQlbqHyGt7oZCou18vrGfJ5p
hgfw48LvG0Vs8ek2/fVATS6FZiJPW3goMvZTHydyQWxfOZArGshbI9nfVBa1bWnYfXx0z9XXFhfL
L6/IyYzYTvPWc2B3g469c0k013KqMK3txDVJsMgo2GoRHeHvnvbamKGY8Fley4jzCn0ijj2oepYE
oBVF4ishPLq4nrrxP5+YZY1BGVGFwDBNpIA4MAG2iWBkTpxz4X8U2T5woigE+BfdWfwMKr2HuXi4
Ks5uLbIwjxXvMglCSzeCWOnkewDGkvEASG2zDl4PyFo5czBIwcpW/pJIANYb71g23eIlxlfr1Sr/
X5s4YVFazzvlXwgGo9UaOyUs+UK9ZBTRFxeu0aZKKWHxQ5NFE1a86Yx/L+gOKGRPqW4j3dCBxXqk
FSgGJ0R8KSdxDZqLgTDMMa41V91k9HPP3kvf6IAmY8bnMgPquPrGkHFTgKEUYvLPXqmKciGnOC7t
d7IgUSUY6c9IzvHDYxKtdbTJeNnwkPDlzKzxf5gybgDYUrsYKbKddmLNLLMpEURD05tRnkrRQiBO
ABgSTv9tcRV8UJJ8cfcdN+7zrMiESMSsU6eFJXXTPrSAufuT/sBGVCbw2p/sx57I8WNBH4/Ku230
C+BFzX113MPhZhkZwDnU4+ja2pQvhNrG8DYVHFUBU2/eCo7KWo4wbWETjEurfb4gceKbDXmhHn6Q
RWRukDGFTSCjlkV9Zd47rBCfXJzHyr+ZFc6jSuFlgrT1mVOXisCVbb1sSbx8LJGLIaJESa7NQMRn
io3LHaUa2mk7cdPj+vFFF2+3ZIjfXaIqPqMrISiEIJWNqwd68OW9rPrAR2MYfrmxMbXJTbvkq+s5
dNFJaHhxHkHiOqvUbVhXsNQ+GIYYIBIEJdblcDcd7JJwV6l0IkdjlGS1yDQNkNLWbY+Ckw4uzQwD
aC3ZPISPyxM7rPF2BfhSZjh8PEI3OkYSG5ooAfB7hkZ5TJUrYyM76+gs0PEl/Ybo7xLz1I1T10UU
atfGmscKEl4QYmvq9BdmsXxVYaE8NVl90a7LYKzB34yhyV/unr9MawcInUIb68bRtce6c+BOoYX3
jQLEcm2J8exO9by+cB2BrRt9QuHZ8XF9HtOKppzVyvyU1uneDC5PRCODmUOUumJdgGdmigJRYWhJ
2fhv0fT973rMA1PtNG4YftCSYhbE91zc9KX1/PRki8zs8cm6xdClCbEo75M2CAO208l0V3gRW6OD
v2GQ2hH7zoV8GPHd8oax5MHvtfAucyG82OZhJ5LZUB8dDX7+GUHVWg3GtQlhiM27bQKnVYogsomV
B8m+Z5xhNEzP7NIN2NDLOLIDgqGbC9tn5BuuBr2Pxf/fSo/0TQ8y/7eE8fNG+GxG4fmHZt+pUFVZ
3JLSuhnObqGISt0tYOhYLmPUdMiKLLQotijOvxfJFm8AJnloBj96HKBELvQy0GHXwszHe9+UJR40
8GfcPkeXrUvxD4Ju5UBktxpWxM9GZSNklC2aAQhJjkdO8CR23//b/b2aL6whWpx+oOffG9A5YD8U
HrNT3TjYC/kg0WSCiLbLXzGx7ILJMjRolJ3K0kmBFMvZcxeYQ7acfmjPOy1l1wSgY468ATG3Wy0p
7QRy2WMTG4vN3pOM9XPVH6D+Yl09WSWs9BdsomW51J8MA4bFCZDAj6dqwS4Y34ll+5MrFxwLHilA
p/R9WxfKWEJDDmnC4u6fXtCjl6bLTbmH353/mEE0KCAz9RaCq0VxFw1IFx+En9nnHMzVnZL+KQTo
hHn4I8pUNyfHomx38xAuOh/MgoN/qMsOf7f5sy5mrHfY8qDIoBnYsnoFTMzexZYnnnDBQnaB/X4u
dfQ1Ei+zDUBy3DE9bJhmbhWOFY6UscwdN9CQDsVodDzfDQRWIWWenQjd6rDHCjFfW6vr3eg6LB+T
xnDh1aqNkkMkPXTlQ2bRzz1yV6jIRT8hUhHweEgrDBvp9+mTlEepDdh59uidk+1ENPktGQg8lOF8
8iTkLIDMJjYLnAtK4CbgIwX/ML0ObtUvTdHB8dVp58LbpZXhXEw9hS5iEOTlflMt8ExfrYV+N/zZ
LlO786+e090jpIwi+STTScTMMjuBgdzFI4hURGnWuJSK7besJuLGtk3dDQ+Ni8MW5CB1xitAXF8J
y8hU06LglLTOwko4ifZpurIM4rhJJ1WkI5Xnb8/hqRO/5rthxL86pOuT+0cEnuU7suAKkJKfg3Lq
mFxdpoD62MDGTXl3nSCBVb58IgavongdYX4Wijs6YIeNnCqi9suFqPkC145MJgN3+oypbJlYk6MO
YhnvoKH0iDw6KTTit91g+wEIDWOe09dNXAWX4y6JFRcoD1tth4tdUlCzAtKIb9b4JsU4FUU6HAfc
QWGYNAoq0ffmF6bw1NY1a08d6soRnUuBuLfkLEn00fmqH12+bJk/t48Q1Zjv5zntpjvsBImOG9rH
3hrLM5GEWtYp/0IpCDKJ393pY7veL6PqBsojVomvQwdZspUAMCmvocwAikjy+AUYf/0uyHrLuqZs
rmLydYqjRrerqcHf90srLYnFfg1Va53ikBr+dq47HjRfhhb/HU4cROpIe9I5iaBVzwtmyQDWZc9r
vcRCh7qMH7gGJ4HkZHVZdESmEA5+eSkt5FksIdo5WE4ugZg+Hj+TFnE4M3frDy2YDlCdaKSHlXfl
fy4x//oYL9w1ttYn1OCW6cgSlKHmkltXGbvroV7kvdZqA3AW2dapTAhveLGLCclLKGAf9nRISYGl
yOzmMHWF8hrSUQj6iNzXeIwBdcVCqCUwKlzcoDbWnk2TveqOOS53gHd0RY8NDz1ok1v11dbgI1Jk
+drGNWBa4ILvbSINW+EU12iH7wSHc6h51M5CarpMAAoHiKfLol7W0v2mWVmk/GBO3W0DKamy/CRr
N1BlR5qc4I1T28QJ+x0EQSIJF6T56caNlMZafc7nnX1kVhf0xhJO6BWnaqbVHbzqy6udSalCMso7
YTNOrNXX3gVsQ8at99eCeQw7pFOReVI0OT2eZIcg3fG4Nl3g8CuFKt2PoqFxnMLjgk7IXmqgnkfU
3MIAMmd8AEy6IN8rpK/EC4pJWH1k7f8M/pHbi/GjU6q+Av927hgYyYagzajGRHcQOmmVzEnIKA1b
ChNdzMGzlsxdQ8TDo+3TE0stb5SdsJAfsqcyafRh3nsUgxmbNOXCRdauRJH3PhP9ihq0C8LE794c
VdvXPaQdreSRQcXERGY+2YaxfUwapGoRvNviinbm0o3JkVW62NO8LC74S0KjseXsEsjUQSCH2d12
hd9nbaVzwfi7NYx4xGHgNIEiocgxVlExxF4BqwV7LARgLg0A/rWy4vq0erz6DCcAQAq+idvSFDde
Ugpd9+D8HVTAYU7cOSoN9+I1kf+JypI/8rYt28QC/u4Jc2tRQoQ1NYTBpOyE564/U8f7HbkmmVh5
j/Jn7C7RK5uaJ8g22Ffc2v392fStlFmWUOqelO2+TIg7LPgOBw40dy1SFoLTFSHDR3zwD6co0U7B
fLm0ybFnXbnD6qmtk55fcCUY0LWX90+n/lxRTp9BflDfOhYVK7vjndk/XRFxY4esmc6yrfXsVt4/
ph1njEW/sdjurEKzlkTYKbnWyrJvQZ7zXPCS4MB2HtDEV/X55W2FOgSHvNn0785jEHv1ohJHeVJ7
7oUyAGzuOxZbVrybtkvYQN+ucLJ5webbilOCD0i/fs7v1dRTNyb3wXuYfhomuwabq0qqs2vqNat6
SYKRCjelTw7Zx2vWyWxXiSHm3QQNxhiUooA6AKHaKxY7DX8PZ29GWgHkf9PThCQVPe+34mI5gIQd
2wIq7JMlsJr0MtY5yhjymJPOlBxwIHxdwblA2XyC2Jt8fz+ye0bu2jgyyFZ8AS85y8D7a0nXRKZQ
AOWmMNyrCmvflg9Q9hASH3hyTBeP2DsbCy0+HhrJBjkVDimE7nFKq4D7tWF5FkJ79GHZjdE2fYhW
Q2cIEdqRtE0gpBhoKilQqly5Jr/2b0M5dEhUem1IPwG70rHxgngLiqsO1+MBDW29q3lSi1hZB94F
YAvQaSVz6XuqyO7Ae/4uxOA7gabrfVrxFWXuqWsIg7u4ki7R7IhekWum44F+4MftkiwjQvwYmND9
EA/jUcW7K9UP7I5YJ6d5DgkNMKqk8dm+HUPNv4Lehhnfie+sP/sdLDqIPobRALMncNv1j2c+zVmx
iwLSm+tt4SxYv3F+zOnmEn12go4bC8Z+WMFVvJfbl8SNBc3oAuKvFwd7/Jb13AGZJ5W9na7NfCiz
oY8FI+GZ3K43djI7fZUcgHZr7kN/6RqU+xXrYZ+xk1r2kyqq9+JkrHwDytO3akOP3hXvK86AG7FY
uKx/QrFuTiSnX/a6d/qRM1GhWfkTMxxvkesobwKLIKZ4mrfWRqNxfLHzUT650gVL2pEk/HQoOrLR
4dxROdykbefreZdpPVq71WYzqb7odbUuPfOaqIdHtdKI0t2LMopCBcpuF+lNmKErNUQtLyj4hiU1
duZf4NqA0ZWSzXj9JYQpwyf9cLa6GTXpkJSKJES5h/+iVYJ3HVaOtu8s8CDW7l+5HsRLTiJSh7on
Nb4genVoAn1FKAsPQA0+tBnA5yRn+ThpLjeJEmRLjo2weBUC5Z7hwBKE6w6iYNVR4qvnvf1wqCgg
/QYSP7lk28kexBeWaW0LkcLZkhYCOJ0Wuqda5fdTE2w3jLpbgA++eQaBrFALOiI49B+azbHdVdAO
+hsGdfBGgC8uTxYOzO8NdpPi5w86TjUmuacdTYg/OrZfppiRREg0RDt09SI5Ijqh12D0kACqHh4T
KbU9A6nRLO8re16fEqDAvZg60RP6G5awt6ESlOnaELHrxiNs8eU9xmSGGE0Ozx0ObuhSpcwB/jCT
ujkbbBQ62zpdj3GOdNQw7MEfitX62j+f1/hLR45bLEapwR/+MxQxulyXfkXaauUCAZ8+M/EzhWdA
/N5QwDpCKJEwU+J2aXkpuHG93Axk9hXEB6Ph0Ojx9AX0RpLXxVTmO99DmlJhmIEZRyEDzYwh3xNb
KUYupF5v9EKG3LiTLNnEIT2QX3Z8NblyTz9U5hWx4AVefEPNKsVwHW+kqrpO+OdRanEJevtnsbKs
Z+pffdh0jTdMT5njGHtRPWhWhEgLXifveM8Fe2iCY/1LfOtyDFpBLcluTSik6UkdwhKe6srIjJlh
v/KPfWIpkpesAwSP3wf1hAIrvdreEj0ULKu1V3q2hA2GxeezvDWAFs+qOvbIh6FWoi8M1M9I4jpV
i+0uJE2h74b7+Cfi33Ff3I3iUEfk8TimiPjjtzrNtxaC3RCj9YO8BKzRFfPcN4S6VqFDJnVGMd2/
rvbr/LHUpQXVCwEhdh2K21AiomR9YcISrPxR6+tPq5wU7z2wvunwRNN4WFOQYwc/IjrsybuAwVd5
6k9gxISyH6FjqjbUe05JQm0auZaU3PI/cPqX20qLvlTsIFrcCXLC6r5NKZMbmhBpdac5xBPRfF0d
e9lTQHoqWFZcJjx32rhyDd2hwlrVh4b5SIMk0yFW4d4pTTYDSXl0JvGb9uCLw+Ql9P4fw6mMhDf5
bfWoe5fsxN6SMUIOSVAoEaikgWYoUdQdg9jQSn3KjkNr8kLuizV6EF3rPCxTqJSZdTVNY6jLTgC0
Ngax/NRLJRz6NSN/qB1VQWtyRLM8gO3IStlW5Yfb5dsIS/ZEPnBs5foIGpTsAVdi+ufgSJWFx+ma
ZZ9jFkbijiqr7xMtjmcBzWVzmwCJhE3/bGt2L9fSzdTEARqEbs0ltfasCRog9lymLNmOY/dfvTCv
j8+5YSD/0+ecwiyVLQQvXOqU02jHZ+AVSIq7rCF2Vr7xxnd0+Vwh5Te+VPxhGbxUSLijqEbznwCM
fFJ5pT+6DunaAhHRK1jbZG0XNQtmm4X84E9kUFeRRYEKZ6nv3sHFUvAhJH1/6+/4NqpONo1Fz5jo
agFdCPjm1ucKV7ew4dhkamEbCE4mPVj/uB1DosSc3d5v33p5ySCB07WMiz9+S+HRHLglTDzdWmta
0XLn3WwwBRnsy0u+fZoda1Erky7uSd59UyYbvqQcWl/KFd2vvhD9rlWCYbSSTEPogZRjdozFXF5u
RG6MOfEwZNAXn2dxajYHUbx0NfCFq6Txst+Kd428EFxZc0ld+81Jk69evESAPEmWsqiNlBO/ajsa
vQqZYCn6wETSll/F51W/PPZOcau8gq2jOKzNJTy1izThpAffWFJxXsMvEfp7APjw4hg0tt8d2tAq
86SNo3FmRxoBUkBwAZjbc+XaBFY7OG3IEia8Wq85jEsKEePCzfrQd03hnKiMRF8swRiqh3WdMXmN
dgiwFcwtTWysRWYBZJFBQ1PiDAdpI+cD2aKVwYwfKE85AQrmgbtLqzE34i8LQBPyh4QXE9rxeS7a
ym1N6YBW4vJxaxQmnmHGs+PPnJWCslffcs5PK+HeiZe1pHBoU3r7Md/12y9/tsFZTWPVxQahk1NP
YCqs1Vl1blrWeYsZjWILAsg5vukB+dszXAc0xcrkP++GlbQJm4QYFsb2FJ8ZX41UBbVBPfDggmW5
wI1ZU8OuPiWj1iyFX/e2w6W+2Nwh4Ya6mnqHLt7Vc6C7S+siBy6rTqYjShz6+AJaYtjNYzhAh45+
rarGiJjf40MNZDyq9O3yFR96SXcUnRbqwGGal68CbNid/6agB1EyspsUgMWjmLoE9H7J70wBN7Eb
Wq9vScDbov9Nuh+oM1Vgk0O2guF8RRt3uHgk6Dgn9g8nAMZpdBCHxDDaJUEtd/cmlA1Cp2ilsGyi
7YpAjp5zXLsJzhJCHA8kCPu3t7vJoWPsOL7fOM5PxHVDBWX25ftrM1m+a4DzslpsumBw+0JIwCml
wdpIDptYANvQiOk/xXDS4kJVwR/YaXEGEjJF7O9Yzjxg/2fstY4APbsw2iIu3W8t2aWbqLIwGR2/
u9J+nGO4sL8Zd0eiAa3+VzxdZiIz0xSJLbb+fQxWR5xCUoR1ySqbsNAMOpqW+KC0VbC9LkFKuMcx
nMJJssHGxowVCfdZFSSao8e/yUqCiy7fB6+YJhr6POHSNXKW+CC6ZEHl/NpPDYCK5rejlWuQsrcn
koaeyHvdRkJ5WSCLf/qBCtFkFR+J5L1xkd3k0Mbq1PCX6SLYbBhg/UEPchW9j82Mjw5nSrODxyE/
zfLiQueZELXmTynuWE8hv9WKXpB/C3gIlgK3CMqHDowvRwr+vsPVRjcnyYRq1udKhhMaiBeYcEZS
3TS4sZYOroH2tjMU9cW6PsKV4SCExOyHUi2mQgZJ9acNIGBCS+1hi3MdgK+gv0UBoZO1d/G/jPiu
Yd4uChgp9D9YMlRTzzniKu26uAZN6z0MBMMME8fx7cmgiUKOaUyuoz42hz8CmZ2iuk7rWwDhwZRP
ak4wW/b0KoEVHaHX7QcjltTwpyWlzfsI0ZnFwHhNhznm61RtID8DFq7MNykZoH+ViZuHiRGh0yCN
0WBqWRE3uEihdcX3Gz7nrTUZZTL4NtoDyaPLecyxdkAFuF4zIotX01C7/sadozWqWDfoGfYPBk8d
To4TMmckFMTHxFO2Oj2CFHk9vbeinThsTJF6MYtt+uLu8318WNsy+R2lWAe8DXRiOWnyUhWnXfYW
oA5U36FUgMr0kM++AWxByaSTc50h8NRO1mU2vMpMOGDkfXLrMrjkVImRiWFSLl39TjUtZWgmdgm6
kocPzo8u/4/5MDklSmnR3VQIblBHME3Qf+Mm7mBoKV8E1WOdJVu6Ub4DBNfBwT+sBULpkqzyKf3l
1cFAYTw8jkq60oxmoNxPNAWKXbUXz83lBWMLvz3cYpZCUX6h42pe/snnsA8eNwWze2T6q8jgsbNS
X44xtG8NnQfJu8hpxNeS6uOfQnQ2PQZaGOr9Mq++lUGtJXxjDNK+T4XPpgcFQL7w1f3E/Jyzv7Xu
B0mKCOqyDMtgurylIAwy0RCFSfPTbfX6uro5cweNIRHge7LgRkbSzxJx1/gbu4Cc8RSoXaXl4Inb
lGwJaQkKvKHsEYd5xw8202OEK9cP8T+kx9i/rL32GFaH9na3rKwz4EA6rLVNni1YkvsORYEp9t03
K3t1Df6PRVmQuk7uGGMvhLID+ms1f/apQeJpaw1ijjrexzMlEG9zl486QO/qF+GstwNgH8oGrXxB
+s6nf4diIIIZAex04ErHi9++0lFwA+uddebtqYe9qOfbYmQleWFDDS2C331Y/hGmRCne05v0W46c
+rsAkfJXT6w29oqNnF1BNoay4/oRzltxr15W0WjCGxZKq6S3qqz0YxBBwkcXI4av6mE/c6uwiHyn
nGglxKQtzDFqUK30uxLvGpTuJy2xpV0PLS2jahR7OovSaXI9dOq5LWj8UvEopCJjOWFvrh/pk0AF
slEFzyvsge1iruIP9j00YbMKAwZVRltL6db1205kpXdpIAX2868iRrfdgFEris3IXOsmPYO+6zTj
5xF1Uq4yHCGm9vJz1yp0BykLJCrCpQOZqeCwkbsHMyxTpacwx16otPQKK8V7q8Xhvnbt3gCoHqP9
bTdxEMhpSTiaDgvLsJCXwGifFLa72xX1+TiWjOsS7liE7uYljNAAf+b7+xz1lytCCES0D4CQQFG1
uKwaTyycBWJ8zGsqArQeKukqGqPp/nKfZRNnbEG2wv7U41420osTGh43H2QLuOAvSxkUImKXUwJb
bryjVRI1h7nZodObA/SUZNUwmnYkXKhXrggbzfqZsaEaLhuN9dJPUwz8DlDFLgT83yb2YhvpLYxW
9ye+nkKteq9+1MCx8nDm2yWoH/EGGz86tyy43IrtXoR8AA7huoftcbqSNRSAqAuv4NHdgK3kqD3N
HnFQ205QABuYS3ISJaCfcGgjXORgrvCE9fcq2W3H0pKWI200dmthrMAP0rpl8Z4i/T9L3gA2tNGd
hanwYp8AF/CfzUZoAVfxBAQMxR23kEOgEUra+rhSFd12I7ReSBp0fkd8YZJPB+g4+M97qw4/vgXV
GpZqlW7r+tR6OEZkZS7qd/71vIJFPKEAtedq5I7JPoeNXRRd7QsSyN3Di9Ab/5Df5+DKXfbV/rl0
sQs6yw90WRXVQ5/GRObHmdKdS4ckWjve+phGjvynAtVbtZBIwJWxt0ubZC5MDtTYSYps3nEcYqg8
6MZvg24oYPeg/cVRdMD5VkSs28O97R5bIFTBvuKvLGSFvEu89+gHsm6WQP4gnhvvQSRvwH397sTu
F00/IP0OQ/zc8MX/tj0zvE+ddKAzLEbAkyOIOFJisNIzeYX1nQKGXF539nJYEntpsmXLbldw11U8
WbKu4fxV7sHMidayx/hrHyLr3Me+TgG8sPJlihPxJN8gaitRwTb0l4f+D5Te3juu15XB+K94PgPV
4/34lSFnjR1nrnQaOKUGLIjI4mABQC0nM3Bn608uwtuJ7PQw4Dsmu3azXUu48eJ13iDnCU5WleGz
JJhsTLHdMAJvDqIJgZvnFbxzW3RyG6g7Q+nVKZfy5PzJYWeB+JK+7Sw1JISjWapIFEIo5BvUlBd4
jbuGhs9Yh5tXQKz0j+cgS0L2+8pesfzu4Sw2HfJN4tJ2TRX61ZHIJrZdKemq5HVYhdHv8VEnbiWB
/KziFymApDKD3WwfMiPqz68SQAHKzMPPI0iSymcC5T5qYzc36q9ubGl9amkdpD4wPo+RtOz1F7fe
9d7MzkcnpKH5aVkDTaHHPHgYh11hDRsKULZiZVd7YtqD+fvQlEKf0AahscwYiPPGkipw28vVbvQX
qbXDaNFFrAZda9HIY6Up0gRe2J/SIvYqGt7QWoY8ii+hNWYplvWkzr4PlwVYG4yVtvlsSdzLACTH
5Hx4G6GkZGpjX0zcYMNfBF3P+JhzOsqPZkUEyVWa8M/WVNUoZOKe09t+UU3GNdFBnZkc/WBR5Wyz
eOYUy6p8FsBjBmNHEkJNX0bpF85+YF3TCtJN6shkFmBpZE6OmDsU7kzdqsP8DrHew3uR7eaxBZNa
juo7bteHUN8h8SnRYSrpaRed8MHwWYgxoKDKDCCRdkY1Yk+qFTUMVaL8Lrl/o7LJJbJ9XbKUrViw
YJhkG4joXHsd/2fCH63EnddNCZdFLeLIzk0O7w7BxitcqZLXOTQDKlIQCfMe35zH8AibAtlz9xsv
yXG0cQ/S++dCuMTK0XbG2Q6mVVob4bug/UqZtPw0uodofDlIcWQ/STTWfoel1mPMxUSnM3w/zmZp
EIYGn3yAmdq5qCfJrAT+2SQSo0l7UC0ErVDRgXH5YemiadRo1WVlM93VZHj67gdiUNl9S032A3Th
xvsly1uc+FmrOgRqd7O7+P9jHaNzuJPCsILthUJEI9TV1u7B5y3jApiNOJIZUiNZ7tuY5u6nmeGd
u1K9sflTxuq1/dIuVe9QG5hrBztlZN193KVtOQahtptwkrm21+7onl9ia5cvfxab/3TZVh/dWsPW
AnyAiDVa9RURbgIXRSptZkLvL9fmhvoScNT1NvDoM+AKk1tf70YB/VnYQMRJV5QjAfiGq1qF4Kwi
VucqONdyJ+l3QU227fXCSRGGJVkH+9LOKm81/IN5FoQaOsr0FzurMDRNBbAoOlBKezBzCG+Dn0Cm
tUnX63hUGJIjXvZtfs7WrweDEg0Vbso48ZqgyV6jHuhWg4erBNOaG/ZenpG3jrgFP2dt5fRrtR8a
BjH8pdDEOGDViHUkpZ90aNtBdXVVys46pQjMzMzh0OkGOs13fCxUgNfquAlMuUeNVVFTaxnzP5ZO
q7wu1rC/P7smOGclCWPZ5kRy5f97lHv3tKwJ5FWY9m2/YUx5ciedmngnQK1BTNfIIex+uikrItcG
FDYCVjGNv0PrplRs3a82jHp++Jw0btkCULnroVo8Od6MJjVtcmBRFhRsfVifJYDCU62ZxLIeqvip
17ZNdCqfulvHm0Pl07asXFg8gt1rxjE8B2fOMZwkNg5/CQORT3T8pwzBf7OZGdrxvOaDtOneEgTI
tUnqxIH8sSlm2Ia9BrUnmXogSdNf5ivUwnEwHiCwhEbGCiYBnvB633hvux40B90ZzCmyocKdrzlX
6vnopDZok0UJKuPZSceziNsrEsLh7Ynp522I1Vz0eNEpMLSYMH3sgOimuhatPbMOhyLhkH8duSTO
mG77f8u9q6aM1lSfO8qw4Jrpt8TiPpIpmTZkE2w1H4WkQcQJ7X/S/1gxIdbtSJjbgxxpacuWXCHo
6g5EAFvE3tmoF+etZXWsjDCdI4YZJogD7rBI0QQNLymv+BlO8E2HUjAbo8zCl3Ma2nEwCGAyR7ye
xBvPQ+8GPWyYMgUZP+YZpej7UBhiWvsTXQiLL7kq9OtmQ7qxVwvQ4n9S5hhtt5kvpshJBPOVjglp
+7FWROjyPtX/98+H68xjQKOITqK7JK1nT8mu7Jpw+17dLjolJKdg4ed51YuoGyHv+2zcmiPmX1be
dre2j+ftUSDDq4jmaSN+GR+iFoA32cZFisUhi96nri/C+NxwQ5m35RX4BZ8+rbtKw5yl9qWWPTfq
FS8zyQTKu4sgaQXvNPf6IFxh5xTDZGSXiTtEGShMZ3RD5evenhnYNsw2iZMrZ0ZiQfuaYMfQDL1l
EGn0Di4Hccg/S3lXftRhycgLY7f40ylmTpj4xYEGa52qPPYXCWbCmuA7bEFRIj2DNwvgPZiTZq8t
gjQ8I2JOcFEN/hNC9KjJSY5HE1oqdqJ4RP/Lt/NdzVm/hoLQVEymF00qJnj6v/Kr4t5hiehVnOp4
77uFumVSWS1PvxQOuaWXZ6IPRqVHjbaBp+hPLY0DtURKEDaKw/wQATegV4+t7QywCVUcWAqMdZjx
3rZelJtqkrnpD7p8RK8QFExILIMOuvWwcwlRvZdwtbxKfSfWoaFhxEMfKiNzwefCSbgAuOld3lSm
Z2ci+pHFCyuY/f0qnSnt4MTLSAukwt6sQktR9tAA52QWJBY89QL2pm71ucYrZmE72meGeoYlqP0e
Og90OU/Mn1L3n7VlJ+I7hToWul6f1KEQvGMpKJAN549tymo93I/7sWUkxwyzj6xFUAmr4q2PTs5U
qXRSvTeGJL0Mwec+dt9IQejOmVaXCuo/UTQ71sJOUBEjcw1HGK0DjuH/KF3gdtAwJJry0yQZnC/n
a4haVlGxq6dFgw/vIaTlER2yaV4MqNJdooD79EgiIkb9XBkmfT+98slQHTNqu5xY/ybWBHJ5dZ20
OJxxj1LlY/0QlyWUv1AShlfN9kJUd4PfKHbljJ1i3pMemXZsTIQ+Zz9UNN1mTxxmByp4T+Tqohu8
UDRyG4z4BUyjFnOgpMFW+6Fah/u1/vlZdWPfbGpvZkc0vW+NS7UrpGF6GGoLeBXDZUBi1ANsN7Zq
/7z6qgEkRBQxLWHe326EG16Og5torcxVoHmIIhsiDWSTJ0gQ1M59FRA1l2nIdCpqBDPRytMWxFt6
iqCXhkvpT+lyn5XiEqrlYKQ6Kmj7As4phFatCg+rxj7tVnCoqMmRuL/pTNYOyRfw7TZ7m1qbyzTq
20jvR+nu8teOwklDf6C3oJDZGxcw8pIg3mGE4GKeej09muLiVY1dvfBeroY+X3nCRP2KYbyhHdj/
F91uvb5W3TXDZcyPg2SkI5a8JCqpkZGtn1zRyqFiIFOIuYIFImQlBiip+zdDPNsYpd8W4QHWW5fg
mu6tZ9hkxJOMflJjeCMWwG/wn4USGiuHBVSTKm5qou90e7jU3a+P3ntHcEeWNxbaZkJhY4MEKz8L
gQHllecT6dr9pw92yqkmo7j0+xx7DgOUCkQPpfiEbWXr6hQTwJN3NWKV9ghbeXMKhZ2ZQja+2Y0+
v1wdsBajTS0uZpiM6cSy5HAdgHrnEtH53Wckae2WJd/dBbhmI1sCfMNxUIVGvfcSzem2p+xXnHUf
y3ekSVyYiLMb4RL6smnQ9jqVDYTnWgCsFqS7/Y4FssGUmuFLH573mywElkUKzHiKIpbfn0mvClzx
iqNmx+oyQnKwJqU7Cst9sv48bFAM5aTIkUTYmp+CKY+HNOsDFb1sOgSZX650QfIZKPe5D/ZAvQp6
GrMtpjliUOqy1tK6/37vUZmjxodROxjshiJiJ/LFpjmu3Wwn/rV+O+3HcOw1XdP0dF9hPXWGP9gi
3gRrDT7yiGPq/8LOuAGwN2nLYTNIRcieQRZ7sNrkG6a/tPk3Qun1ib8A0eNMAEuNyi3Djibmw5/G
XVC6T6v5FMeYKnsDyirUfNnLHgdxjdv4lzzfCl3FYZVIH2N4zCknZeP+vLFBP/99mTvwrWhwzaeW
zLk7Y6AgAQcVHWEwe4MvHAft2hn16ZK0y0D7LJ1VsV17v0cMFalrDo1AAorwKBy3PW7fQwOhczmS
gKDfkEVU8zKt+nOcCgPwts9mTpUr+8UjPAMghcy2LqHoszICAfnYEJEr7VxwRvdJtXMYQ+Y/95bx
ahVRhBJvV+nm/fCUXp1ZEU7VuXg721P+BP/EAKg1VrYzDtsN0GAVsKgfvufTHZMchdtfuhLsoMv/
It+QiYMJJ6MD6PsZvX+v5+SxaeoxfZTWArcFokNz/FGvgdigoYoDJiJAoSShLq3WbwXxCJX1UgU3
kIKPzBW0Wat8B4F1bG6/I0V0WTXHr/7nt+K1SvB2hagByWmTllvS3/y7xhYtx/ca+Imk7oXsIOkh
IXTn44XJ6mQblW/Qk6e4lr7+elZ6XpadriaR3iqrwheNpeIyfvnuCVw/GKLj443p4s4vbEkSnt8Y
IJz6/Nc7IKg08L/YTpXQI/aGJ0o3x22h05jM2a2ZcEMBXSOf6JDSPk+SqAgf2dsGZZp62pIJtDRc
LAy4Pe5UeMunkpm+dcBXbsdw5/ooV3xFdZ+kf0s5IsTa3q7uoilKAeFlQCxU9N5u2R2ohS21Bt4B
zp+DMfJ2gMT8I6Pl7fwoE/kqPGfJybHSo6C2qiAmEdc6tF2jwQfIty52N2Q1MVA/kyXnAPiRuMKZ
0XQBBH0/vqJ7fEM+lFhaTaWIdJnjv7hgEnL7C1cHZNsEFza1O3FN/qvs+l1S2baJPFiT3muUKbz5
z/iSN23MP1sIQLmUIOLJkTMyWRtdhASNeQWWWMNNuQActsjcBELkBs00U6t6//iss9qeI+WxGlFG
5UUZQeQFQdkNqn55QsRyT3pRPeGA99SNKjMJJUFwSZuJEnEzPnGUQvgSsSZt/Oq906Uu8m16Chhd
xG3vgkDxwxHe7X54HUHDRtckNShY/cMMpbwzU2g18gvXB66DJTluFMsD4n6wrNqVlk3UU1cCGtn0
0enGtnYBdYJQcSHsRgRYnril/rVa5O40+4XyWjtane8/a8KMeGHEbWWF8nbM4WwqoXZJHLjqgi6b
AMYm0evNk+5zBoammleGEvQLhLYtYKINKOob6bYfLkoups4+XUwGs0MkVzF/NuE88tH8v1RrQNfH
6h4d7MynN6lR8Jo5/XxbqUzc2WSxugp4IHgMR6BUVkeVuW2vpRv7Ded11lxPmH5Sr5CQA38f1hu7
Y2UJRi8ifpzETyOf9gZcNqzlviPD5uoR4yP2X2M8JwVf1GjlZjrFAmAa+ynfWmvw8Ii9G+C7+t2A
/XhnoJtboFmpR6ssdDjCP1SUN+sD+iMfRTkzIghJVYa7KJbF03sYmD2byTPiOFSUjO6s8TWTlSX9
YYX1crJ1W3lmIH4NJF/5S1VgXVz8ElEaNsIVEdbvbqgKegJedUiflexlwiPhuULI/2aMWSPGRfqf
dg0h5u8UQCxPZS2yilb0F8rzLn9+oZVS1TkCLlrBGCruKASWM5fySSy4Nch/rOjGYEjzUM7f/wMC
kg81WkqpvoY3M0kHFqjV4Xj6iVp3cVITOy7JHacVsbg+sSdwe8scboNAIMaqHEmtOLPdJ6AwIRFr
kWWK4ZnclgJCoqmfxZh6nHOJMMyAhLpfTv6uxo5OqKUbjXi/OqUthPrlYgUwIRegRcAW9k9ctpCt
dmywTAnwObq47OPNNtTvKQVGbJBeerQ/VVHlygqCzGkzUCyv/h1Zv9LSe7nIJWCEJ9E6VkAdrSEa
1uFkmYrwQpSCJWn5K6ObVPbscohScucdg5TXyf8B7T7SteijXbX/4UWXJJZMX/HJCerdSvXZB7nI
p1gua73+fAHV7MjGwgN0jFsobvE21kJ2bfZ+WzS8jv5+aZTzGNB+kIu167xE6qAipssEvQJagCm/
t0s5L9+c8JDQ2eVz+aFVkGnfH50Auwc7VjRqLv0wljOr1z01srzaerK1NnLlzhg3ZfIRRH3kq8Bf
+Q1HmTrc+MEVoceRfuMElm6BGl9bJJa/KFDzG+t/qbm5FeYf7KAZl14rMdLKRBFgpuct/WpkVl/J
v7F//+5MWNLgM2BVOsT917j0wTD7Gfrrg4m76Rapbgd30o11EePskiCJ7/lsHRqY6gxY5QH//wRG
6wg/SaNObct707H1BLEJAldge9QLk5anGu9mtGcyuNXf4MNbyZgE/Y4tt9PlaBqjBai7gSoomHlA
7qdpR9DDOLdpOwnkqYDBcSxLmCmuTBAcGIpL8CPhBYjvpxYE2HVygJ9Lp7H8b61rE+m9AFx9OjlI
YGRB/8xXin24jEQmbEP5ZcNnljR9ejoOvqVMv57wGaGN2PKHm4IlV+MDk6XOdKpEgJC3y0CaVF3r
1IH7OiHNlGxmCP3r0E0mpkGM3+znRBYC+/oSoZ/bsrAJ6N0RRdGXu96Y6tfYoum0q4MlvIHCqeXx
oDVJsHE+BurEl3Xwy9PUoH4JV6MwT/QG5Gc+qt6M0S02MGv9fGnuustS8vLu7N0amslPCQecgXll
dgoIxrkZmlJLRdlT4fMfzOV6hCa1ZrlRsLOdSGIW1VMa2+CNQAJYK7MIuOCOiKReINtXBGA/w8O4
dgJB8SueG3yvHhKc0PtUUao2CNCr22yASLJ7TCxuy+UdjwUepup65gcxwWynL3XaEm+QDYLlKxDq
ZrJHBm5IhwfJc4hX64bcHiTGC9hQc4ay3HvURKOmDxrP6tehIJnPDzwLMNlVvLL/fnDCPEZw3i68
nRG+57NpuPXm1Kt7Rd2ArIGtAJ2msxkfu8heOi4rsEx0XLWDVKLqlEectftp5EbabT+SCTcvO4mo
FfMf4i3WsK/cB4fAJeB6TX4eNiJmKopDQ+n04PX/70bfCcANWTRZLRxl2EeI4/alEM3KJn+zt4QI
4pO5x6fQxPBOGBQ2gJqOzG72Ph4NRJzhDxb2As4M7Cy8Yj4lRHYZAxaoavcHyaXt0uJgcsUaKhyU
TAhLZ98sS+bHW92uDmMmDQHxSMM3/5lLn1v/psXZnKR0wRoTCGX1Bv/57kuBYutmYZXyWkILDzj5
tRrG120145dV5i5tjJsuM868PILJPeXM2PYdJDmhWynB8e+7+EYm7c60kch4E4lzUl20wumRIoNV
GQ+CCmLPLjBzJybX+eba0ISdFjJLrugyUWHwcO7/vScW4o23byeNADrWeu2duLN8tGEC+9tlYnt7
s2GttpziPImvWD+VqdAgnUkfby0sFPp/CMIA7vPK6W8czkvoV+z9eJ4YY3CzmWZtIWJPVw8ylhh8
im0omxM48CdFvw9qpHOvG/3Apu0o33naZJWphzcQI2joNz6Qd3cKt90papaahTgqXzUs4jKFdpAr
HG3djWXBJGt72Kv0Ii+4noT9E7J3R4w4LqAJaGH3yT+uQBCQEKbkmxlaB7GVIQZaIhzYbni6KKFd
yAnVoRHLG6WUpm9Edv8EfDrTMXfUphVIoSalnmS9aqIz2z1m3Fnp76Lqm9lP4qGTdqHOXFYCIAwb
k0sQy6dyOlxzDfmMtJg9GNKWm3YFjKgyH4ZacWOEF6yxiKn7prJ1EdZOMAj5bfLctIlXoyLpltKV
BHjJSwEukTOx0+tsSiuh/k6/lMG5dZW1fkCB3ZkdxkchzgMtsMp54pR3Qz2ZuJtRk6iOeEUzUmA5
oC2pfnGkj0L/vLMQn6WQr0zRUMcPUdFnavMlzprhXDKyqoTqu19R1nMxm63Z07HXLPBV7yuzAm+n
X2BdHxwPgSZbHdrejfURB9AwCcFaUbnJL9ONyydlZ7r+3odHRZ23YMoHsnKY+dLYC3WMsgC9BMXZ
MXxHpREgZXDafJxqY892JcF1wdEW1MccxpF935ZSOdVGw4PcOT8yBikdIwLId70fXdeSbocTb3Ud
DYnSpugtAS1NQ9oo9eDLIg7ipdwfZ0xovIEOR9ctzCXsbMlIyroK+wiSoDhlJO5b8IhfguQTgXmB
Nk8TFJy71NOEOYJKSKiL0VkFZ6NCzVSSpZFwVRpylYOmMu0sPaj8EuLzTung+zuwBulkptaZ2MJX
X6RZtGFHX6stQGiOEskAAMMnHxo+FretOYZpgHzMehMvb4mr0BG9UE5NxU0bossn47oxbrPuO+JG
RKhw+Q4DoTMG997FnwmJukhS531ekFi4L3xxawO7CXYrKKA8JsKA2WqWtOfUnek7PtKD10XUAn87
CpREfufJQg1ZlwhgwoYFEAsGKOwahgEgfidygX7bd/f15De8rZGGAvPmok+Lojxr9ehLPf+StJ81
mm2opRfC6q1GE52F265GeMpS06Bar89+URpAZPDvZvkgmRZqKQRbOrnOaqx96/itFaQxxclEhfRL
aOu8WHZqn8/eFjagPr67P33lLgv0KssbE7i0dk+C46vBh/diXdKbRCx1X7gJLN0HIhJvE4NMpvVI
xzIF4udv2PL40DXb+/biv/MuSMQZIZ0cJ+K5Zwbi5/BR2aB7/dt/7+93RBCpUQYHgaFTFcx2LBp2
r26oGb8upGWmjTfdP49CsIW5QZtZ20VS9UnN/ZGffdrfl+lPzYZdqmGhJFHlh4U7e/ip06kMq98+
ZTcX2zvcP+FfXyiVBzCreyXBwZn2GjNUg0/kV5+prLPV5/XyEZrxMV0FMXz+FhbF42/SbYwbzGpH
GpIjVOTJkiECtagrTW2/NXomN+2ECqgt9+lLl9aXqrbSYJryLBwAOBLXn/OAs3EMuWjlrHwlIWIK
M64tFhc0ivXo0U/NqHMaQjUYXFn/NWKV2PJOSWgfvpAe7Ai/BGNrBgEI7/4ATWXUaMjatoxo/AYa
+0jI7K1Ngk3PNnZfqGV65BrAVwdmywMHetM7lMUYB/L4oe/tDPKxxGf2pRNLes7yWhDJas5R9eZx
LEJUEYg5C7wFY3DAmLygg3VSEHY+SJytTQr3uUktS3oiTOfQjw5n9XNRJ2bmhIO3QwQyucOTX0w/
gjKfXLcpLSMaX4VSexgEG7tMScfs8FgHD3AKSIMzJ7T15kqhmJc4hEJc0Dj38w+Vn1ekg9NYoN4j
sXmlBGhvzeylDg57+5oWHlBiJM5W75HE8xG0yu6iNUlnLKApLVv7lH272SA8INHk6fjQavJQp+mS
suV1EkNfyceOeTKoAj+MfGm4BNgX1lTUqHw2/8t7haBoDQdY5T3wNozrEWoIPcU4GYhae6Tvi3qx
goUhbo3F2JndQDvUasNQwmEXmREhkf7Zc3QyiDdV6b8SQGkuo8oL1PYb9KxZ7PvhAGl1nvPO9lgj
WP707wnQEf35mzfHDPm2F1sshpz2VagTk5OkNpnjej7gogqWesfuIZUgdtgdJBzUdQgR6xJxDIEt
Dd16sRJaDrDOry1jj756lSs9KVdK4FxCPRbIzvmc87/IEMFnE4DZSL3okCa4XQo7NlxFAgHquqv2
Fn79OPhaRRXTlDIXcJPwR4yItJD1o4NZk7YBlewhpzL08Rw0I7uXaJ5+Ut/YIOoraYyAZWQ3lK69
3Tg4YMM+4xyPCQ9Y72GSWCn/SCblUBOvjVyl8pmNO/7JO37VBe1UZLev9Yl7yK+ouzC84mp1y/Y4
bQEXC4qIdy9wDLotPVWTlOPgUYxuNrmm5ABvDVUBuFPOdp2cc910JY9axoFmih0Nbnx2vLFq7/ig
jzl2+UxiwOnmbGXWiTYCQXC72lejXh8fJpcJeeIOelPDRAyEy6h/8I/xN7l6elFz+6QiD7Kkcwuu
eNFFSQGM+VyL+GdYnpWes1IHkTc/ZMqWJa13WcbOQP5TkHYPDt5wujWC0aa0NpWVdO4ayWNHTo/+
yvVwLVsZzjRKCTSw5YRZqHqLEYpm5PUbwqLfvS967IQoh4MK9GKo3gTOnW6xluCMitCPWcsv4WE9
fRoohpWEQUd0TkCPaWpqme5sn1803BbVpFa1fHC3RsKv7cdEKEWb06epTYj0PQBxuO9mpQSbiQlk
sMt5fHkuPjb6gANlk30OnjLSJU4LhwLHVeVf6+m0j+xbTnVT3oss514+2t/HpDzUvYMj7o+QVGT2
nIdNPOIPHclItbTuG1ITl2/amlE35fN+8zFTNWez9j4tE5cdr6UdOClrJ7V/kdfDieo5AyQllIZR
aqA2BUCguB/rBkhkS4G3wVxxqv1tybZP2jtu05s3clw5U/iRx07Me3YYc/PgD8vpRloU3oX+J9DJ
mdQJlsOXQJ9ANXefUCebxdkIJtmQ4aDEHlv3A5wag05ISN+r0d1vzfhuE0/paPDQvqb7OSeeTzYk
YKbWzNDhnCuDmkhRy/AO2+OBxV+km8ofFg+nZKqueIbXoYntS7zNwUDMBbcSLc+fImW/fP1K5KiJ
ad/V63QbG8R04nm/2gpCZcp81nVOaw936kZeQ60ohhfxCdVWCbQWj9O50MVrGuwQ/XAR+ruS24nH
yJqpt5R3z2sJ8ZeiJiTOsshfzPSqjLkQ8af5sUxlzjlkXwN2VTB9AlcYr3BB5eVWGrqrpiCdXZ+J
jGftAoEL4PYyPeE3Kq0nGvJsfnc82/I2crn7wz4JMwhUnl89EmTAFcH2lgMbaM391KPYd+gDrMRL
1Hry7VO+itpMVwWruxI6ziRQpX9KV6pQcfB1ouMsKuef+K3GBofa5UEs7lUYYN4P9kDeyw3qeLHS
7sBD2mk8yAIGNbNs8kn/vbYL4rnGT5Wj/Mo6/fCJcEHVJuNCu8hYymmHAjhlqdmzblbiYfg46CcH
JgU3UI1Bd8hAm69/TeruMLPD2BcsyPpmyictIcJ71Mcci7/Q6aQrH6rLF7P5P1XZOQQwsbZs1YWj
S8nPCqMorUnvZ5KPHOKiQHRknY0xnHlQ7lQpQM/kNkF2rzduRsPETWTfGL581qSWhlo1D7ezBGET
a46kZN45YzYsSCLDn6TNo2+b/7x19vRfHr3SoqLcDKWT7OU8VpwnZ6Zs662vNQSQUg9OJmCjMLOL
Srr+rSSVZmDc/Li7AD7Yq1NeZaqoiF8X9Tl3/4QmJn+Xw8I9TuIIX5bTBpfNBLceGC7WW0mNvEUG
nX0MCGat/0Xe1DknKb1JmGoWIM7h6fqyOMQ39FxZYYwM0RybyR5evhKBwbTz73erqG951QlIBT9D
CYPo2guV+XTu3DAkIaJTmMyfgqZeV8HzMUrDlA+t3uE2p94KPxPfHESGXsfQudgww2kNl7Uwkk2P
ig3JhZ10J0apE/3kaqx/qrC3Php+VaHsSDcuqfqfeO+KQGe1ZO5J72B0k81r6j+q3MkgE3ptkmQE
JOI9PzCXSTzGBogft6eI1Jppc3LPjNioAn+9ijCEUecPjhP59CIOegFhNkVvfIoAd1fr8go7pEAU
V8vy0GaVaTmDUlQqa8rQgq3mWrmGCD6vzvFNiMOTuWwU5x9razCFimWnW7WfDK42U7Q+k3irumUe
6emXyCrC43OXWCJbAVEAEPp7EHl9tejSbXMoiSKLD6WjjC6UptMFftsopOQQoE4g954O9xosUcsr
tGxYVjGSX5o4ojgAiGqlk73Ch4qOwFJQCIR+eJlJEAkzwp08susacvA7VPCaWneYkWAsseUryBoZ
50z1xrBKrcTSXkxQQlskxA5OdeDLK/BvWfXD1B59xhfNMnUu13/CQVOzS2qEI3bCOSCe9ZJYWde6
6cwVtLcOC9B0gR9SwQlsLQZoSTHI4SyZYCXFF8wCQTRaxcZZ9DDwcVQxBmv0PM2mQ2tDCjPGtMp9
o0vwkwvI3VgtrXINgxEZsqkPzhhFcaK6G6ek0x1JOszVXFE+6AlmlLsV9OJyHKVXm0X2JyUVC49Q
QS/imRkXyIPbMHab24yIdjanuS3K6qfVo3yhWbDVwBREnHelu1HyZOrzrhyVP0DJdd7GMAvPSNa4
xJcOW4XDR1vajonVMc8GAWmiWtek+OzHBM358velibvZ97uaTiQToqOsBMRw8TY2l2fW1t1+3MMF
PYipy+Vn08SU93oXh6q6ORmh+ztvT+KqqN9e7OOHa3cveAjYib60YKxJvOFlKfYH9ystxU7s7zLS
eTsCuMobLBvyle9cp284Z0I86JSp8mcOAYN1hNw6WJ0NL+4C/krKcWMWN7Y84EyM9kQF4b8cJxam
LLYklsj2tLT22N3JILl1aKL1xWX1TqOBSZ+2tKBJppz3LhU/HU3cvA0P5COrPAuGEIfZMrE1V9Xr
7dI5e6ntILmC/iBbMtbXfVy3HnrOpSjVO/vJ7aXpj67riGuYnvdXEcMczGqIFHNSNwfHBzgik9IL
xe9Zl7kERfXcgrwfWAsoSCaJYsjr2SH2RFlEg2vTBi1nFU7ZWSd7/hsKnVz/FmTCq9seWymQLvrO
FJh1DD29kNfO7KuioBVLPkklR2ID8yVJBMaEDpMZItVPds04ZDqCKAdW/0x1VeWwXs4A5ET813Nx
MSaGfPLdukvNmJwvbR7F8pXxTx2uRj5urUsqDGPfbvEgSbwIZcQTTZV01Dj2EeawGQuSi+KF4xyk
Xl/tUZNnXvxsNyBTdSIiwHNGOhiMweNh+Luc93nsknAERFICIU3cbtbAdNCm8DIwgUEEpQqcEUeq
9991I5lm+E0SGoFTHXQRjOfRBZzjQoDxltuiePtyLb22bxsekThEwR7bGWK0WdliLp8vQfePdNVI
trstFKOoneNU7YYFeIQw94fQEj3myxbd656hqNSWthooZb2KCEpuU7FXpWE9a/2ank1mzQBaDb3o
pZyt6qhSNGipHOpsnDLqVUiwZl7hOiAFeZ6cevGMNKk9mG1UlGUKdrSAG0oivxji+wBChS8nSq1U
bq736XAWG5ZelObcVa4x05ZZcPPg4amFxfCgcX9R0iS7EKt4gktGgalfE1uILi9lqfsOSuAeajlX
4d2KZmWf4cPbZIlGTNP9ELwplGOw123SqZcWFi/x+0n2YHzrXfq26wWBcXOWuq3U3/AEmzK2Isam
t2OjaI8AoRt46SFPs1veGDYDxHCjwFXEIcF7Mn1usb+mMLZJTtk2KEq2H3M9yV03rpufXVeHPBoW
O3Bd7Msgxb3l9S8ouMC4Ch8PMDmSJCS9quqaLwUjN8bRPr7r+BBsm6ga39Ur0D6VMcoU3PBxPc4P
SBuL/0nSby9yrGcldIvn8oUGCmr2KQZGs23YHrllurTW1KN2kq8eHszv6K9wE3SBaNhI4p8KTT0y
egpJZ7n9FLjZUnHaSbkbTSmvQoQyWegUYS3ewSdk2AXuGZ4z6il4/NbJnV1r+zGpmuZ9oZa7dn0W
NpUZfE/pvbrBkWsDAOXzq2DRtyLSl1ClBm1CMzhsdFRFVheAIYYxGBR7w/JaamA8M9TRKwM67Pjs
/og97nI5jZhQ0Vy5GM8DU15sJjDdE5mQAGIjpCrdPNP2mJvseSBXVm1CCfI5cZRkZ+pX6hGeCzhz
5ZNThR77PogIFegtYuhhdgM3AX10QAQL27hJiRofftGWa/EWqG1aYN2Uln80jqTejJ8SdEIrlznO
bzAnlPPOBszGwjDogkPDmDC8tfb36/r6cJr5GcQJmEJrV3j8gwk4OF9UAzGASrrCKab4hdH6KaqX
uvNA2N2Hn9CWd6+Q0fmPfIeRZPgyMsEW7nMCR4KIir4dzeg4gAoTV8XWSBkL5sWMGrh1RX+ZVE+C
rZvwi0pfIeQijq9YYLCZXe6B2okT4xmhBKDWu6K/sHKU1C+kG8U9BAc+XeVvy1kMAn9WCpm+uIFC
71M5RNpe7v4zP8ft794bNstqrnTMNtyU2aGu1S4UhFSZtWF1w6YiFtaBPuLjvgndXJsP28rdOi/8
J3GgTGsMqf3FT368u4syDd7J2iGXwsGnGrcVERoFLefjXle0zTxTjXZuUvEoyBVzGf4hDoLAA+Po
xj+NQ9XGTFTm5+rZmw7WK8eGWAk3OJEqVgrPUMOE33NoqM5ZT3gPxL1DJ1fkZH1raC/Ic1p8v5BJ
4chbbZGazzLWKFE1ysWh8m3+HPdyZLsWGX+LyXnIUF8PzfukZfgLZEE9qBGqJxwqh/wcOPn0TZN/
5G9fcEYL73uAUVYz5Z/i/L9ukqL2pfcujLjVaKe+wuQZYwz5dXcViZ6KuASpCFgwYqkGRmXXXKDS
h0Sb3MhLwwM14RE0FqfWlZgSy1WkvbudAS1FDBBlZ26xzRNQtT5DtNz0yiILb/VMInSZOJ3ypJvO
/C3bOSi2DVqWYHqt0u5EMkRfKWJr5nKoNnlxb0jnItraEgddYu8w8K4h2Ae1Pi7QI+z8TltHQPz3
9/giY/wCGWdX8amYwMWkFYE2Nj2gJetnaeLHK3cqulkjiU4CS3hG3hMawKVsll563HW8A3ZLPck6
DS0Xgi77nil499usIpPPoJJQWiQmfJ/1Z/8Vs/DMJRkPmkiaWAOijKd29vuqa6hs4MPmwF5KGv4q
oiAjHavkEjeuNveUfSLtzVGLEmg5EuiSkYTb0vicmYyDyxzScMO9Q5JoZMJHtXuS/p/8zTXrmNQT
qfnwYY50SQu0horc/INuFnMeZ0FIkFhHCKXEPhZw7xHW/fU18YslSAOHRIXgrf7zMWMrmdAthM8C
EMFWEahZbj/Ta78ZKRusyuAycHA6hSsJfQjfDzIXojptrVGkv3rVKNMeAa8EpOZeQQ0v/ayzw+F+
1ud0PQwsAYnMiM9Ha4CmIWV53xQlcU1H06j3rBIdbx24wLkh4sCQQHV7uGfQL2Nsg26zSgUsiUoY
i4MKvnymQ7kDAoxR2LWFj8n9iy478nIQKdLPWVG372r1UZjUyqGKu3iV7Y6f/1mf49pAIAxZHwZY
0UD2mEZJSiSEa0Gb1WFR6Ht+v0ZuEf5W3fAKHuO4ql5T/QGDWy6OK068xCWk968Y2+3uod6kpeRi
F/V+F+PR6HcZrIgME5ftr2d5RLRNgeoCukmLniQfF+/Oe7Pd1PQtAfUT3cemeMupfPLnzYWYAxFk
2PqBH5IgHXcuguW4ngr9/tLcsJ28JYcBeg7JAenHe4THuX/Q0MaeFJVluWMWriQSi1GENMXjTN4u
XYPdg4r5CABqp9fFL29bLsHd5APXHWrI5nB7N3m1P1CySQ0K0h91JEEx/pBg8Q575Of4scc7YhOE
NNoFdonIOcNICmFk8FgkJvuAmuJPKz/pThZdMTW1WaOeqPibz1z/FYZtR7XE8/ZpEX2lereqSaE7
yEkxDAXjtEya5hqIay0Ioy2B0/NfDj/0wnKrtttLdrJVZ2pBk7JZaMl5frMZnQkR1annz+FEYP57
ysT7gk6i93hcres4X03txY6ozCQgeJNSa8IEIhcQT4PVpCV6hr4JA7XcqsBzmQULhC/KgGco3LHD
eIAIRTvp7DT05VZvGnouw4tVdoedd86mKVRKyAszNeINtnWhxPNrgFg/rya1w5mZ8F5P6+6kBPrh
FP+hqSMdXYTk48EX6UM+/UFj33oKrx+ZIk/2EEEoU9dWQPkhvSuoMDXzYnmucPjEV3SUHvZHTEQR
tUdS0k/gxqRD8itllWhdqbFNsofOqtAiehsGPZ/sbW4lwUR32/jK9YW+QKhODGWbTyli3a5zvkFW
AKFU2TsqR3apONeCx5UuXoOBR7474I2H23NOLNKn/xpNBuxdosJGKYz4beMTgiiNs15+q1f0CZAS
4EJO8CEsQcgNf5dFSjDLQ4+uZyyHDBOD9k2OMImBL7dAMTDTRS1xseLwtGSdQzB2alWVgqclVE/T
Amq7zVdl7Gby6c6j3AL8dcd1cQLhATZMDX2YHxI797gZ7j3c2xdDwSW0QgY8aagFXdtNq84Bm4wt
apcj2sHRJa5nJ3lnJnqte1tSbH7ND/Osd0MmgrIJOKbuE/+ksVAomt1MZYqxblFOLaalTQt2M5va
oXGHvu0o3jXUmpR5Oy/jV+2AN7m/QKbSHdFCLHfiJ2PI7/6cmGietnT8ppeicIYYxp7fYIatI8es
VVrk4X0Y79mbdPTYoR06IZJhvhkiEYMFDmKLiuqNBzB/q9roBhQTiqrAar/ZR+Ojfm2lKyfTNvlc
B1cjXhsP2J2oCXifQ7YFmvZrLfeBKbev740ExmYIhiHpn7emdtvLzLB9m8ZCspQWznoRchP39ZfB
oc49vSoo7ABE7Jf36NS7e+Vi8Iasqc30loB696W18kI87MfY818K4LkQ1w+Z1tqIbqWjoK7lgAbw
oG3s0CeQBC8C8BR5bKAHjzC57rV8q9Hw9W9DqxtDFhjkOy9vMO27FnOq0smrFRXV4pRz9+yhALnp
JA0UJ52bD85dQv13tXkUKCnlRcB9WY46Q0ynTDf+ydn0dMHCfCV5LgU1HTN+nwq1USFg1pw8xn1w
/tpBRMVUHOy428XBBViM/S+SKbbOeUExJql4w653+QvYULgiNOt6Q30hUXKQh1aislSyuXSC36Ho
lXiN5S/qwSt/YmtBvi6WHWKvR/41asDu2YvXQi9Wbj07hNhXdnJxc5fez/0FOItFBLIyyraWMFH4
Xj8m/GR5QRY+5t+sOjJXjGIk0JoqiYNhiD8a8SAIYqE6Mhb8GeR1T3F8mf5h0VOmEGTEaUypu4Mc
nD5Y4HUDBwHULj5RcjX1TXz8x/tpoCwxtvj40wnK15J3qPlMYZd54V7/snrjMfODHMfY1nlaL1tM
cVt6FsUWdR6QURJMFTALh0r3cg6jSyQ2QBIKp4xKPPr3C0y7dT+fFt9BaurEW96y48snzi+B7+Pk
4OK66uUAp/mMRPPWT/18BTstJWrtOVTmv/Ze96IGrFI2wJrV5q9JrcMv8qMCcLy2e5lNbdDwEH2E
pwSYjn82UR1xihlSGsfTSXDmKVzH5ZXKFcCknMLS2LV5Tmnx7ezceYJl5m0yxODL02svlzoGu8lJ
QU/T21+gYs4gGR2YVR/+vo2qxixG5yoy4/OqKO5zlFC+z8UD3fsK/Z8CBtEAMcIy6LfsesU6j3ka
4w4b7tfz3xjWX83uuM8CR2TTZzdS4LjeZ3cbNShdd5OJ7j2nQFfOD7+Bn/B+Gp4bb/tEu4rhWBA4
RCDBMPexDduoAz6bgNcJb5HIWVK5Pk9405bisDaQoAE3/32NtRqiTCikMO3txEqsx1XHrdN68kUZ
j4eoeMzlyBpG9iOI5oKhQjxpWbTlmI25l1NGrL5rOW5ur/cxhScQlepTEDxLTe3TeXfdKahiAmDO
yTBKreE4sK6IdeBY2HdpFGVQtiNBmiRe5o8FTc/xlrdTfKTPNGBjlamBOb269gESJGKY0oe6vEEc
2yU0tRkAOJKHuPNLjYPIc1L4cbdfP05kK6rIsp2NkjZzVvqCKidjbtZN3VtQAjOrzM9uVFo6wNJx
Y3rfG5p0UIRsc1T+28vrzM+0vqo56TDXgKmHx0McpbjP7+PouJ8LjL6d9PrIV+azbDDpnOcz2bPo
eKWisAK9lH5jM2p5/bsl3WfpskrIMIxgXx3JrdiDKpwUNtnq6+CPuLzJSL6Q/LRdytRR8AQMb3fU
8Bv322XIxyPzQytlYxfu+v+0gE4GW//gxyJfuhTugajfzn9gKaekSjNU6L+BWBgEHtavYldggFid
0OfedIGxy09cRsayxbEuvIljTRb8ZzGzpr9qK5yHWqw0KZY5XTkFiTmsouFOgls4/OGr6CWLIpUY
Fzubv2DWzYk7YN6zqAgV+WHrRuDABdAFTSYms+Q2jfbzUX67kdiDIMBc5t7Ari5qxrPR5ZXTT1CO
Crv9iwcedOgh3cFetGeOTbpSUJrTvnzWr7lKY8Ftx14lxWwxA29+7eaVuFwswvERtapXuZFgVYUJ
7JDqdAyGfOV7ldQnfq4nsBsznL1sE/ayKFT8IizTYhV10KtHPjM9BPtUTlog76eFDMkm94mqM5r/
C5Od5R8ywo4T7PnsGsuugPMg1OgBatgzXPkvHFstvKMv+fqkLAi/+eD3Y/j2N0FL3mdJrfS62f6h
ROBQmWUzVXOvEoiXciGO9ZpxXwdz0gufGhDfAdGJqr3DTUN2gwCbVv+F6gRRF3qToigeqecXxGbJ
/euNeh0FfCpOY56/UpLXhH5ogCrYF8ZapWtNBCKkcFiGUxJAbMkOAEOXM4PeViSX4IUJau/8Rx6k
Y2XXfkSXKcLBcfMB/Qa8AILgS4QKRlgxlqj5x1ZqEAj11S5G9d6/n6St0sm4GdffkImjaD6lhcP0
ClanG2lJIhWrL4r7tln4u1lryojtYT19wIHMukS2BoL7apfI7R3XbT2YHSvkPYalnxFb9jMoeQkR
WUQ7JX8/8DoBFKHgMf8iyABJxk5PBUWHF/dxn4BA7NJo9eQWed0pPqROr0vgW6btuG7o0sm+CtGQ
vpVSnjwbynDz8u1uXOnYosoC/0rtwA0t+nqw/4Q3D2rZ1/ynejZ2T7gOGSuD2VIJNqPFiSz6AiVc
/UK2sFXCzezTdYABgjo/2WMVRarbyDo9sQeNl4Zs4Ztmpy0z4meB/eLwV8F6iluhEBohQMANIhAf
eX0SCKiYkCrdD1LnickYlkkIgFwNrgVH6J7iHaxatrIl541EjbfAJStQaPIUZ08urh0r/tH5BOtp
ruqw3M5xNwKGv7Hzcsf5EX7A0pDKI/Q+Td2YsetQdpZSFr7btAtIYROxJdjRDHFj/ho1tgdsD+9H
7omQshCsqiKKVENEvKSk1742I0g/tZENfv5cCah2toUS+XPGiTrUVM+TxZVaUWzoEMhg3BSEuTzo
NwwoNpGKm1HqwwoYbp0YX/Yw2gzNjYYYT/9S/YQWiXTDUKx25ZJHdsfsn7zOC72zU9Qjf11HX2bq
rU+yvdbNB3hdNmaVGw9LYt9wWLHfWExxalX2IJjUbf+u2Pv8OwwBYb2ID8tp6xadapLasJF25d67
rb9ivojYXS/tx88udSn2Xf6J+bJrZrln264DJ6UJcvlEPongPwB7L663nNPJce0B8UbARfFQM9Lm
icWUXWLNfoYKVK3OU3h4cjEYuewcGee227ArKBQoCPj40QJNzsu8vJIxLSNocxWU39omzQ+KGjA5
sYg3U+JCMKeZxkZm5ho90dnQ9LVRxZR3Wz4Dr3Db//IlgLtHYUjtgvuiaTB6liC3Y1W8lIGn4ACS
qgUs/mcAi3tLjfkzI2AwQf9gbnoAYSDb7HZaapGHk8mw/nxjt50QAcCLPurBEpn4ZXmIS1gmngtn
VLIL7QPeN99Y0S1/n3bhzggz3Lil8kqQj7nuhIGXjM7Kfvw4I/QCjT/GcviwbkusOun4LsQJtM6V
8rxFdgi2efzRVVdpY7NPA/iFyNxel1duOBRQdJ7jEaQf1X2Ig918zX/H1uaJVGq4KDf3WMd4YBTM
nu8l6lzWVRxPf/5/XRJFcE5vKFlyltI40A9mJAuAvaABX/X7DuAqAvd9EG8W3S3u3EL50PGHl2c1
YryjOSsFm9G87P7ZjTjrO7Ak9jHHJEzPJBNREgVtpPmeiISYkGW+2dEr6suoZ8cTCQo7WAJYjr7T
rSw+maWD1S/b+KmbVbJdAiNpmZs9QsYd8Ni9yQVZ4/2+Vd90478Wq0aqdAUhJ1/ilXdi7UxQl/X9
Gu9XK+6j6czj2gdF48uWMyhSfGabCn1e/8YBuPM659JVggFPzFhq6UGdSPOCZ/qL42em5rcpzfOW
DbPTNOfUchdNuaDBmuRiv+1dX8kxuv5cs8SFeSFQj9/oukNEn5l7GL1eZwpG5qO/EzXjTDWI247w
u7AYd4NomISg1X2P+McZS+2QtYqkYUGmoEeHaYCcuTDyUSc4BIbqZ+asmlOfkzNCgXeVEgwDFXp3
U7GlPHDLvN7n6yNQFXlvOAu4REB1auN/2TaYRDogQMCDXRClFfLg7BzjCyd1268kevwjoBiKNcKD
R4J8znwPS8r7/PfEDB1HYK6qwd0GeyFYQO4A+4hhpxYFku6Cc++zjCjnBWq/t3WL2vJtkFaLsJeu
h1DqVPbAg611V32Y270tiJTmuy/jTDrd+2CsdRsM9/cnpTUxQF43WO3ltdnRedfJVvrdHZKveaHD
MzYZqP5KPeJ+8STq16yjFNVB6hOUPt+PtC8F/Sf9ijV2Lr1WjMAdLtfr0sYr4g/ZqHStC3uaKvUK
iPeBbATpOm/tv72Y5kEou9oFfYafYYq7oLE0lCVRPwK6oo65tb+nCVGWh43GPOJ6wmuiXj8clvFq
nn3dHNBz549+/boMoJOHRHkZyi3xjFlnMDfQO9c+ktMiG3bqeyiMJKx4t7mC+CX2HOGrRDHO+NTo
wObse+NX2onhs4BxsyUa/0mEiSqajvxDI5hzYDF1TBc9FZcXu+PiibKxuUz+y1xzqsDuD+gJAGv/
5V6rq7Cq7Y10stGnTc6b/2yJfljeM/if2mPgwakkq/hj80G9/cGyXCrS9jQp6iyKOxqlzAXaJDei
o9dvwqyHTUCGyrBAsudf84Sj6LIBMhqVL0duBR9rH7/ioUM/7TFG0+wRk9WgNmEHeAqVGs+KE53C
+ryeQvlx12/5yNxcPR7k9rFoyoORC0FGvRu/puna5pI4df/Z78+LRpVFSDkFV+6TMHnKTBrQN2uB
JOKSIJLvXcHQCJQyXkUcEo1LH4GKmmgLs/+NH/je5e+UEuqBHp6Rx2AWFuh28n6L/ahJVPp4NROb
piE0LGtl8Zsdx4R9UsnBFBksI2Y3XJw8Bv9iT8tjEjzwZcKrg6eJI8zC8cSQ66JYtUEaOjHC7V+V
5OOx6H6uOZg2ZTIKDMmXA7Wdg7RPaM0ib7XCuvCsyHuaSSC4lVfk7j3ApLBK72Ulr3ABqZzU++5h
uBJtEJxSPMrS3YHZ0dBVEDKSUDKDN0pvk6urZaGuxbNj0qpjulmRN0uxTdSowPxU2tcqnRBUCwdv
vzc/3ROXuoiBaYtWWgzkJdKZa1I9nx4Vh77QGc++0s6AtxBdyOMe/jt3IHfpvO1Qwsq1bHwbY5Lt
CaseTZ7cQlCIfD1x2WhmlUuLr8mqOkeOLgnwaU3iycicetHO2MH2v02k8wd9X7p6IInpHrFMJX29
Q2iHYcb8ASGfFBMw3I3Ao++Bl/pcOtVL2YM2AB9RqnspD0NPCIXVuJlayVY6Vh1gnkeQw6heO4Da
0pxwstRTuricxzz+McOW0Bjhqsq2wIBE25Z40Rr+2gTqYkidAM8b5CgVyIDtdo22/Wg3MCJyczuZ
q9alG1JCWT2h3kLl22AK/8uqJHhUUB+9vi7bZ3VOqXZdeiYIOHyudgiI/ZqByWLolJPUvwGNGtOV
zf2yCJZe/GuCF47dVyqvz0eQ01cH1boICBrcEEEaUZRb4F4So5xh4Dd8Mdoc7uzf2i3Dklq3UwlP
JbaVXslvcdwe0FuuWuanyInX0OiELNexRS/sy/uNgaHTd24Th3JYexm2VYzkYbHaj5Ee63kve+oP
wtWpu2XLj53sllvrsmnsVLc2lQ90Y6GBOPEXxCrlEWMJcJQJD0TLypWD7+OolBDmbzeo3l8xpP9i
UKAy76w5caRm7sXiY3KB23qgXGu3r8lLTEJLjU20u8zDpt2L7v5RR8LUEyUCnB+Dvl7pWjTL1M1I
/84bHQCQP3NAuhOD4ebWDYPNvHQko8vd5GB9ykkhJ5N1C+Abyr0FlXq95WpqlXuQKO72FnaR15oo
Z7qlus+A61oAMLQrCQzqT+Ja/VD8kfZt9TaPb9AqGZP1+dK9QUqJIQYMjzP/v4afbHjIUFqA7p46
8PnfhYpRjEMm+XsI+wes3kk2+7yA41naT1daM6/Ht1Etgr38WrXzbzN/1BDIHG4nBgRoxOmPrNZE
RIVYkvJowtRpc28Ay0/7h4YiqIx3fOWvua5YLFjgyiUcAmuKmyPi2668ouzE7KSVIrRYXrjkEWLf
WIytzvvcgFcgElMBJswm4e7mcERvmJmDHR7yhUiZ98EnJAIOb5MIfXWH8lerDFcCcWKR+fRLkREF
7PoUHLsvjIk/66HbhCcUw8WqN/8wFXQ1qqvGkQSSfQrnBmoAXi74R5RktsvXmRDH09RoswAjV8wn
ZIU1VQWguzI39JoR0wQbgzyzog0bDMEQczdspHXmzyiUPeopXMfShNUjVhjVPHqiLp8cPv8ZH/sL
a3xiZcVFb1zJgcYV9tyNse5DRRhgakMQgIpzVNpxaTtLyXdKlBQoULz/E5UX/bgSdodx0sIpM0/N
EV8WtwoZjBZ5Ie7C9k4YT8HCsZop31ECMfxrnqck+NCRgUpsIQNwwpkEWIN8z2BbRDx+OHJ6vQPF
q6TtQE/f2i3ARXSL2TGrnYQ6LIwmauetXNz4D3qNTdJX4G0Zl1+mMl6ODoDiu48UIivFS777xc9C
JTGbPW1BOq//ayGO5IjgGwL5LYNyjPHMep1QWGIPAVU73vAc95Hn6QsdIGhSvJGsmqzle+08YAX1
rLBa+eJc9aKpEvjicT2FUJ2Is97TYS2eR8BbtFXVJg/aywXHqr+1rD4URl8uu5QKWeMSCRVPFBvw
9qfLTtOm134NGpsuO2M0XyaOe+/t8ybuevn+kehlhAFb9PkKEwf/QT7ogNqeD20Cqwj8qfux4QhN
Q8+hgkdeWWlER/i7WS6kLwI/XIoDhd67dluql0tbJhAyQOuiFsfkNZk/FhoJYLh6y7Zd2Lg4J1xn
QpSszzwvcd1kZvvXefJhW+Xk/N/tRaRp98Ua9IhQsByalaGzZ5BaPrWQkq+PLfgkRoEGtP33jBCu
GGhHTGhfqKtjx/PXomMQ22kqX59/lsiIWZktmGspm/sMU0mP4JM8YVqu1FFn++v+kf1hkgjfAloT
4fSIdrLLEONnpVBdVRiLIFdFXmAqSe+9aVS6vVz+vbf9szA9O9fsto9lk1rzPllUwK1hPwPC2e97
EJ3lZ8Pg8yluyRZ/T/yvQYnQ4Y2bTOpPY8XRdvDMQF9iX5pNsDppuPgyzgvfta+rcNlV3IaFBOTd
f0KXcDsRk7MCi+9+zB6HIP+0TU8TD6UTNxzKRgsic5lRTy2lykXApPhZ3Ni6hNqlns3RIYEAnAs1
GdMbH+DfopFKzxmT04dyatl/8a1mbkI4+gy5WNGXY7veockTmXpxBqe/P2V5u3Nl2ldqYLJm5MsN
6c8KMuTjfZ16Bfn0wDb+j2Yp/t3l0R6Q3saQUPbpug81l8wFhPKEcfV7IFWojIka3hotoDgu2bO/
zwSLaLhTgTSJeG0OjYGPvITUq/lo9WUu1VT8sFKi4stzvcshseSNAH6Kb+LYzn4gyW0Z7MQyLFPw
l6NGMUsGzfLb1XtW1RKYb9J3c5a/A5xDkZFG5qCg7mUrtyl1IYxagCCPPpY17GbgYXAahcWKGGJ6
yhTvOKRfbk3fZpC8ow3N0AEfW+VZLCUEY8d4GPguAvoXlZJWpAN3kzLhuSY/0OdCz9TUBgIeL7ys
s58vqFaPbfvYTvQGa7q96+UUAFrw5ngui/4JEa5DEtxHLNhMvNujfQeJq0Z/xtyHfQee6kQp6Fy4
Zd7zcTJhGQ+Pm+fsDKqboKUEtvhHFUpp6KH0/HgZA3th7IAUxr6zs9V30k+jqVxz/jNpVRVWqM55
DShJVggme2UZQ9WDCrlScxwCmUU6kFoHtQ3hd7pr75v/Mnw01x+1ur8hJVetOg1EYnMRVwIl1OHT
3s/8M8E65qtW2LsVdwOpFAmbu+0W8DVzjE5XqTDtdq5cAPbc7ziXSP4uHxJLY+BIUXAaeZpDMGR/
SwB5AWwgd4Redc2AyFBI5lM12vSpeRStNExr9Y/Ba6z6yk9vN2rH7mN2ZNKDCx69F1WH2SpkiU5d
aWpXyjoW63zJbni6XzyWgWUjlwSbHkWfXIozybez7Gpz2IhlOOZkA4ArmMvGiRf4GvOzeZnjZgSt
iV846btzWS0tcYnm+PO2PWJfOJCqo8FL+SMv+EcoEvURchWJ78EQkj6kTl6atXq8DVLHaV28wjgw
AqUFaKugkPDc0cqZF85/DY2G5qBQnZlE5nvrxbA23+YwEb7A7KanoeV37TqbUZ94tCnjoMbAvTDB
Baw/cYXwMkm0m2Dcwh5UthFgdw5IBTAKXBtrtnD0cStG9jXjwldHT30hvSI8qpir1ZPalcNGg31p
LHZ6Ale6KfdGfYO/oEH6n2kGl1u4OBIHcMrx7HMR4HmDY5DoTkzxX/e0kBdJnJV2XbhCW4Or+pXt
gSBymTqHFELEltBEHTe1AJYpbvvB2L6OqoSIjxEEt2QUiTGHk/rmfvsJd2/BO0x54zjOhblcIIGK
gVRLoipDYDeQqPGGmK98oF0P3qjT3KqQvtmyKfr5pxc5JD3DEVFdl0Tko6wrtGegq7HO78+C/lJm
SR4MOkAKx2kK0/G9wzSAeNrKStrryUzbM8Aerc7iT0QuxUqzz0R8OECbdh4GXdbO5y8bYe1J7Hy2
TkDglP9K5Rw7SFcj+bM8CWH0UzgwmvBa7ZFTo3CGn9fpxYQbeV5x3r8qFdnFdWlHspcvCIBz1GH9
HMFCD8tlCLYEy/ZiDTBvpGludWzN9uvRrU4cEvZHavGiwGDeiWf92g4oxfFB1B2p8helmG2IEe5b
V4xi2RAl1P/oDz9LJIHLi+gTFwPVegrQgYDIsRumzNTBmtt6bmCkpDwIzKea7pfWZyXpGQGK8zwo
cLVdt1AxghR2giGMZMW6KAg0Nw77Xbu/n7YPG6aLla5ptw+wsJb8VaUQJz27klHm/ZcRZ1iGEyKO
PH3u9DXUdSxdyvaSK6RSf45KNbDic/1mPd5IsEeIIlcCOwE1vmK4L793wAJqGEHjj1xpRl0mjlz9
VQiUfM5PXTfB2FIDi0vgthnuRImH2Ujar+sreT0TLzOTE64AnwsGbXXXLtxq6cXLCoV1pIA207+i
mLnOMoomPMI3jejnB7xmit5guAcWSEC+t8lxflLWhuzOoQK1MpqQ88nKInlFjCi2dQJP0PWpooST
DzjUQCIel2xm0qhjnXgx05/BDKU+1QmRHqf/KHJyP43hHEOrvcY1WVhYoI0RrhEF7AIr+HO840zN
sLA6DSPIgzrd6Lcl+gMwpvxSL9OzhKfYEGXNoaXADQT5zNSkoSW5qyQXyCB/64U3sUwmyBJKELry
YLjb8dv5SEU8EmWKU7xGQB5KCGWkyYI0+oD6UawVz04d8LjzfTq0Z13QCcEy7OvP1lbpW8/qZu8x
oHGmMFZQSanWsADMsWmDYq/ksRstX1xqLWoOjAWaK0pxNdyQOqN0kr7fR3V/YgJyXus8ElpuqEd2
sd5Bo15YxI2oQBeYnMBxcxUffaN3z43cL4dbOgKV+ftU7JdzUEwaRSZ20Y08KkjEZoX3739O6TAj
gtHL/F30Y+GDDqanTitJe3i/lCZ1zaOsMIQPmIyBZNQ08SqAzCbSOhMzVDaesPLgwHggl0QeZSAy
6rOd39VulLg2usgLPgoT2UwFM+DE3xFIuBxdVko4hsn0vC/gZR/6pcYOO9Lfbx7rb7hTHHdIf6vJ
t+3G5Zy9HmqySomMrtOxHx6fLpW7FObi9J5KUZzicQFDfI294NdTiee2mS1q65hiyndNKXFd/Ex7
CZUdoGcXomP7UpF/FViEDejW33x+i+t5smsu+VIqOkHJjCU8rkmfQ8eLjp9dxeK9mjZ/gIKB4UrW
EMUImS7fe9sH704nUjyd1kLxJS6uH2Sw9lmFNWFV51j+Hh3r7VKi1PYNI9PLxLbGEPAFVAuJkq9Q
Q5AuywAMUQo72v0N+iZCPyw2GU8Oo+EKC8NJ6AF0pZpsFSQyqj9GJ4UAae5wZU1rulIXtD0y99/s
GbKc6bnbxunOW94tGCJqHkrd9HMGKaxKc+dNzPYU5Me3nuQZr1UoMv9wn/MD2oprIRVgrMm77n4X
JMEbboUxyasXSkDizlkLN/J9WIqVt4oLASkUD/pAbon964ntSIQNGlP1vgDcPvtL4AXVZhy/F9V4
WtMXXrv+j8+wWTEaqKbWd92OkZ6bvIaQp38+ccG/8+ziItbQ2VsOGHaxXridfJ50CO3HJJOOjEJp
3cXiJXrxhIt+Z9IM4x8jsUj1GkdeXPuw4n91ENsWc5Cf0gGt2eK/3I+/1zVW3Qip9QQWyi4EBvfT
BReSac3IVTtxRBB+ObxaZ84AFhxB0Twy03kuD6qvP+dePLNNuLRu4nuU4a1iGkKsr2MRImuxbXoO
2xLkPIRuDmCl76pZMz30UYJeVgEjh/VFPDdU6tleRaTHP80UqEpRtsN8NDE9l5rGAQXoJYTM8Tlh
SqBSh7kSTfqfbICbUxgDkW5iwW1+1cUmuTeqzfEFIwrWR1EE3Xs/tS7qw5V79bZ3ArbfYa++jfdw
lmp28cdKI6bcORh6SKcEhduYoSFAIFpIBahST6a838jVjqlGgKi08CtiWl2ZjaZyyip6Vka+fmqv
sC1reJ9l1H+UZTP1L0frQjo6UCXAxleF7L+ed2abXT1S3GmZnbe+yc9SdymGWHpnA/HAQM64LXTM
bjEaHFepIvyb21ltHtrDteX+JiGieIsewoBBYtr7clyUzn12V6iQBWXm1lCk40UFPJpw8iIczZK6
/qqEHkT0dzNca6eGSUy0T8kD3vbo08P9o4GuVdGrB07NnvUFqRb5pR2ol3dpF3D9bNjLUymZTf38
KlEzYi2tQbz+W16CnWD2UBSoYQW2/ZDVKa0a77jxYKx0hClU4A6R52oUU2ic+D+Y4hy1Dn1c9M63
hRpJWNFiGzuY1kYg2JKAy0OC+IKcbJh4B/mKoABvmBlpEqpKu7UCdgCCo88TuBDjKTdYOm3GnYI5
94cgcKRzHQOwM90zR9Ujjqpy6KPacVAFNoRiDKjAAgNNHj0hf2Wh8EIeqbf6BJazIRecZiE6OQxn
iA3rJVd+cAUVWeHCeJXZ+ha1otTlMDZ0RsoLJSMMRYxyibU4aZZ2Z9JX9A0l2GHimbriamSKHJfL
keo3v0pcP69DNGC4AJrDztURch9KbHqMA6uyQnSd/GNx+xFzkmc8hDnNMwkg4LzKVosCNxkZmbWd
B7XwWjxgYYeycABVng5n6uviOUnekjk2a7iTxopFrDYhh3XRAOeqIV/iPrF5LrB2ArfgVZcq4xfQ
XCu7K6OcXLfHzhg4wtoSoWTN1tuOHYi4/CpXJ4diBwdJBKUPV6EbX8qhF/9AtUIdlfRE90/W3SQy
vhVjilUArAPceQ6Jzg5GvhDK0B6pwqLNmIZPn0hgazmIb9Y501yXRK6Ewr8KjKirk2kEOUkNStAp
y1ex2opS3OrBFqK+fajMQA+b1+P0oemaekUbgp29JVp2xBtVjnWVK351G+dyB29KrrnTV0wShqxq
AYVjlO44lvNaYE6Ub97qDZsVit2SGLgyKvW7IkmJMDJ4Q2e/rkgkpm4UB29kdLna48LJZPmg7PyA
Q9FmIOuU0cMsifRYIwwpBPeBC5tBkda8RFDA91UWtlVR9I8LgQM9X7J6GX5PFEDpTKpDDcbZZ83G
5Z8T+xkESNX234txm5/gLZuLM+zJ5sJMbGOV6wEgduB5ZcVG8zfbcpgWBwu5iTcLcCy+Im3WuR3q
ziA+1/6Bh91F6cHxnwpWPHr5VNrumg9OXvR5F7/ynhP0/2gUdNR7Wg5y+PvQGx/YSlyterLihexk
xCVU+ERImJPTPCRDAsfM0AZsobhUq7zoQJKaUzPyNyoN+zADBq5Q5lGZrPpk2hWGCL8kgbvv2qH8
maLz5Dpidgl0Fr//+Jy4M2RRKR5ZUIDAiLGjOeLq3YdmU8+Bo6x5bkntNlVj8nF8e3vJilZfI4Pg
x19WJE1pvV9TFmYAqbxJsJpXjCFOwe3lC9BeO3S85eYoXGdkgBJ1vGzQagcqmCdC7GPIvPK8ex5E
GlFwhpzcXE+NCLhDjWx8UlKL8ePBGrVgK0E8/sr+ZLAHrKG9yUiB30OV3asciihWnQ9gcyzXO92F
0gq+mw51eO0TWE54O3RRghNaXjPxEW1zAUkPkjevzGMQf8hZ7L4egD6fK7tgo1EQ7KPsRI5IRnie
+NSJGfgP0qUqkglBRNvFs8AWOu746fuPIBSqE17xkbJSYgVWWzmuyVUo8kk+DdLFYbuTsr47T64q
tvMf+wUdauN6n53dWTRaUb0npiLSChrmxsTTH4osPQ9xKYA1VWqIYUh8vSuAEggFpJQIq+pXHouh
81vx1laabRXNz5qzopSLH3R9c/YjyV2YlxkdbQ7ot39+fTO4gszbgGyilOhGskL5tT6hVEOMa3OQ
Xb8dAQId4GrKyM4PQcIo6uBR0OSy+6Sc3gHgPCDV/h5sxQNt9T7mH+25cMEsjl23DeAhdxYiWRq5
xrYrDbqjMSNax5gffVOGMLpWJfv/mh5atIcdj9S8XSpanHMySyopc0Ptckr8xGEVsBNxL2ETB0KF
4srUBFzw0WY4cHd/16FE07ucsUkf7g9t2gNpf4d8WDGl+8mJAoO2tXKZN5EV1Y7aNFkVk6GDV0AG
nrczkE+MvsuomU7jmGizsNiac+gj0xz6RDTAEkIh8UmT1JZarGau8v0Jg1K89AjJc18Hihw/RU71
bHMk6XCrGm0ND6jfC6FimolESiNJ1mKPB8EFgUH0w/qqbwnC1ax2zF69Tm+2TxThSnFXetnR0pC0
+bFpoPXxYcj6MqhXpy5EmYbmsQBd1l3J0SShEm6ZpiOq2YzRtxgzTWLQ3nUIipifU7dc3OVVkP8p
CuzXzjwnKnS2ds/0DIBjoYM5jagMNq7Colra2SrpmPJPkBqJAxmt18+mK5bBZum6rBzeejxIl3U7
60SLno7nUsg/6c6hONPR2MO0PJooeg4YSXM7EWcWHrjnj3y8ruz9QhUDjDK36i7WfR8fz1Xhyt+3
2k845fJWPyevqnD3H60BBZ/U+XUGEt2WhtdcAUOnIXj1D9OUq36XC/tvuqeyFrg2nnGGeh0O5lOG
13mwa2RuLdB+51CWU40YTbeyN+k3KVir2nKzKx1Bs+UQ6FEZ5wAl35G6l3v20W35JV/C4qUDIyC/
r5/0rZs9Extk9aShRwq3d0BBEliN90vKM7z58dWwEkSMkRdSAliGzJMIKtEefuzN/6dYkgeqq48/
kjj4AMvDVu4yjk0YzheaB6/4IAQvFyc6k+QXSbmMdqmx6SdpIjjDa4+cUZTde4glHVmYFZi5OzMa
oDwuX2Q0BMBS3RZh2Ox9Ki8mYLmO7aOKzdwZcS+Nd2EnfHyqRca8ZG7zQNBjPS82Nd9uVXvqswaX
6imCBv/crKysJkCbegkyYBuwOORDqIN+ckm6uR+QWq+AqiqjEZaWm7eBB83leFaknyFsR6oPyUeb
6JTIRr/JMgY05J0SmjmoPJWFWZRmVaSibA+nP0sCriUtEWEDoRzHCs0E8qA2rxgvImisRPAKyJkP
F4O27KCh2qaTfgGTNhGl+9LKX32AIPsgHXCG2eRaOwLQNMbqZCBJBCpTxuXehB9D/clTo9fE9uBD
DqdqKgibRDGpGXbWU9M2fimt7X4EhltoUHZ470bdCYnp8AslMGZF88knpveKjtijEXKAvZCgurrh
CZ1PbGhdIw9V8mSwj6tY1CBhimfgkDyGAgs0hoP6UT/F30rej54Khkin1CSlNmLnudHvuhcKlHJC
nVVOupPnxTWP4KQIRDvo7sXlswrH82SqGtLyRfNQBVxlLhkxFtjNyVdWEVZDp54Rnhbfhxc7Ont0
JqwCDNvPGtY3N4apuJQVB2HegHHql2YMKFLS18S553hcHlWcPMmoAtW6SqI42WqHk/9dVe+01v1A
KXMS4SG+uVe5iaYSUJfs6JCjQ4DKDZ5jnvXpekQP+4cXwHc5wIPtCwV/CuU637lbdqvq9dE5sC4h
W8/K6ePIrA3FmxKIlO6rbUradXO81846CuVV04L0O8Ob0+2/XHHhtOLKDi0lpVAl9VvmErsVIFmO
NR+JZ/hQehh1GaJt/obb+KjNfEB4QcZpBiRk5+VJ0Z+1wSuR89ZsNk9ZwS+BPQJl1yl+gbQS3Irj
Cp9UmXLE/y5pYwB9MJlLYSbYpNol1HZ4LVCOtCIkn241R7ma12JKgJuZcVM9DdbLBHqsh9jfDfbb
kLzbcz5f7FFLe4/OOsY59xeYlmsylI056Ivm6vNNhvSRDP2KRYujzbv+dgvCRorPAXr0ZYGgkt8U
6oy5QAODIDBdIvNTP/Oafq42o9ixX+hp1MDaPDRm2PuXImgoVVXkoLUMFvW/wlpSFEmw3TxUP9TJ
tJP0UaDh8//TzyI93rvKXPsy2JmjKznAWDmHi6CNLAYpSyrZMXcD//5O8LxkiInSNLjI+cJ0lOWJ
YAvo+xgCle6oelh5ED5QTLK4pnfsX0TvGgZReUBOU54yevEgMMn5Imh/e3u7kyYptR5acZG8+6oH
xEkx39P4/c13ETNNHdk2XA6uG06s0jo/y/KF1/uovWYq3MqDRO7GcZEXrGBlNz6hmcKPjIaTPYyu
FYo5c8vRdR7c4eLN0+whuhDK2YsNz/nu511B92GXUPwSyRLdP0bUE47qjcLQygvH9iXya2tpS0Mu
c50orGwbye3yWgRVrvDQGbz8L126aSYVXwwF86+h6uZrOOaqnl7lIU/ZtobmDP+R5iQVoQEitsHe
rc7PoqZ4FN84h+dyHt5VC19IYoVTtD937GezAtQ5COJbDz4RCKnpamcjkIdOUIvALSgzR7Q4fLO4
EHPtQS2WYxo0GJUF9P8rnUBt0zqaPdwcstaLeIxIXNemlOrE3MNIN5OAkJEaNwuQgDKEOz4U+WT0
wCI9VvD+w8yn9f9NHD45CPHr4qzZAxtuXFzDIIEwOnhdGEvr7whsSh3NVQkw1kTr01vCJdB6jjMi
vZ9h1vHpVQFJ7XpqUPpeBB5zVWvsEUPYZ2xcNOk6BVjvUnXIb9cb/pYaaGB7EjDUATIY5jZQfaxG
Gl4enRjwnZrCvfKG+2t+vbZ+MP0iD6tCthhJz5J0mBpo2xrvypD/H8PAHe/Gu+6mE4E2ARkJCURt
MvPebE4ZN4DIB9TrRa5A9IVh2P64h4d+H0WKpyZzto63tjt5hQAmyhjTiarx80qXS3WYnFzIAY7o
PKnnHrGvXtP3uxREZtJjQJqDVJtLUQXoVdlPUYRDOP01sy7M/+3y+/gUmE20my+6fRRhqRSCya3Z
KEkSo4RhV0QFSgiRQZNbKx9KV6cstayR8w6Um4Cu8E6b4U5xNprkjNvUhCm1FcqQdsggyySWUBxR
1mjiBmFf3rOdegiwE2E0GLN1HKLkliFNLDySJKhMhG4aOhL4xW1jCJcP/39eSFvoPtO7LsWMyFul
A4ty504SZqDjQpvxSomH3Yf+EPr3C2KenMDtuEnCB1JDspZHyvVDIxmQ8sV1NeflIqZc2C65xZxA
TxhbIwWk+Yz0W/ppj5EwvyKBjdt+R2L5xVv2QIkzGFvVmXwZk5jvuvkuejnVwocswa5Ip7OS4WRp
OY3kUqpUAnvo/+Dw3qOJvmcZ860hn4wWRf68UaIrywOOVT6NdD2nxurWkwnFOo8zCIYmQ0Uv/JR4
4ALzEyHMgxH6SDQQrvWQdhTp4ha2Yw0qGmE/jPxpK6/dVk8JJuBR9FqGrVQK/3d+YjWVg6ngaSY5
Z1dbe0mFjPpCZs7KHFVdsM8rcku0WwlcHxus2Tc3MQoQfn4cLHC/ohYtZ4T3VGGPI+Ud/hypyEKl
cr9tQxNa59NaFdoRKdHi4h7TC/qCYC9N/rjVIvE9AecGG+c35wxsetiTbTEm/Mr1GKSkkzZ64Oeh
07OnN2SaIo+/53hHRa6RfugJ/8hwlz8fDxvKuWFGzm/2K5Rx7/+450eG1Ze6R8P3Eo/dtULsdEpF
5bqXDA9qZrpwiQR7/vbcKq4+2BEw4OPh6JuW4PzgruAbQ9MqWH+XgwG8oQiTrKx/fwAxrm2EVJ8O
LiRuc+SU8rMwVoeM+ZQ5zk7XqFErWhthV3IbqVlGjZjeoQjOQpwK3LYV8dyD+1EB7Q821V8Ba0bi
MH0ZA+4+PzB2fQuhTB7TBTytIYATzNdFHt0VsDUZsjJQVV7jGF97C4TLH/05MnbXDqKpmuVDr8l1
7Jysd2dSjwg0gK9ZY4vo++tFNotcabMBgQGEbS5efey7BY0KX+PbvoCWC8OxMim8bdOQj/CI4s21
UvnNpIV3KNtq3IotVasNjkOSYjYiTdPuOyyV+Vx5BPdykxrRmMeoSQm4HHxkwD6eMsfdV3iPEwzq
k4geVB9i+SiJHNVWkqxIJfLMfHZKs9tXE0Za4tNF78fyq32cdKiTAJQwsChCXMqisGLR3+zU+6ev
f8Qe0G05740IcZ3Ng2X+pBmPJJVBFjqEC41BaBkYTKSXOID4k+jPjPCvVnK0mOrpmPbp4ilIMipD
az+jGGGveNmLLOk7kHQzMPjGVBL6n6qHRUx7gIS2x67qK9BEmaBaDl4QMOMasGZMOl52P5hK8jaQ
gMentTtg4BXJQWIzfg17nO65JcOm4uYKBSWgXN/DlyvfxlbnYEs+87YNWPa/yq/Pizj3FWdfeluM
JzbbBtd6Nah1lm57mWqd+ZcMAjah4TrIaxtUvs3CV7hYT3dU66uVc5veVtdDqYLi9SzKb4ZZaZuQ
uHsIpO7lWivKMZ3TX1j65zLLlzCN9ehyFOqhhuBCgJdLT6vNy/uG8+SyUqHIzl0jfSkL/1m3J6rW
Mm5Z9xkDEpWHkIDmsR4E2OeEaQXAq5Zat26UfshuZjb6mt2vCIq1WqAZ++2Q67QOnR4ESQH/Padk
7nCTizqq+GVk9YrZHZ+4v/Gjuw/JDtdOWmv4wBH58SkRQuI0DxHzFgmVrqUZPdCTrNwoeHDt9w/z
x5Npg1TgUHrSO2gpcYw9hVxqUxkr1+DuHgDseu7rAuUZRwdpUOVaeePgtG6JFzNVGrd6V0VpdBBI
vHSAv8DK5ESXOeJtWAJ+1EIsu7+6jcyiAOUNywSP2KpkEtWyBqJvn4DK0TJ+kN8cmzlt+j34n7Mn
ioLgBrlA9bZzmVunQW03iuxTFiRAO1BWNgKLyi56A31W5E2t6ByVNRzN72+i/lLnNN5dKzQuiUJX
KcynNm/evmnNSN7cOcHQfENjtyss/0Z382KIMKsuCEYFMMickPAC4PF08j5DdYJ1DLGEsNGbtNFF
GtFvq9PTlo6xxKlOwoQ6+Iv4eGYC7GlL38xJLMq0zKijg1yzcKDTwhBc3UID9dquIK3E8dH2Imh1
OUn81AvKi+48j36xkiwRutdQb48cGxt7hAWsil3/0N54Gv//peFkWCz/sgVYFFglyFKhh2yEM1N1
nZSisUi/hsXclD6hXIgLKytLYRxXVsHFvNHISMzdEgzjRudqUGYwAT8fL0lKETa23sDFS2sRNXYo
hzuvojB07lo8LFrRvtjHOg9sH+tj6hp7eqwnavYbJ5hlHZsoC2ulI5waCM3qH+jECRb81PCLlLov
00F9uIACuMUeE0iNwGO+tzuNZ2W3h9LAqDo1RHfSOPuSAHuHGsayoVqFFBiTjaX6Q/FKaDhhx7tI
9yxpxoJ1QAQAk6X4Tg5FQn74YNrLN81EjRKrZs/WNY4zh4ZA4y8hrufFqB9qFpGxVRa9nbeH+3mb
jx8wYJfarVIul1nAYTABGe3VwqMx75WjZsrUZ0qrAcZHK1eHfLRLtMEOW+PgVVM3zVYbQddgnduD
CnVFZhsSSUU6ko4z8k6gFd/Xlgk3llNoq4Xvzuy7mRFWZNk06mK6HsU2TVZU4c693XzvN85efPsX
DMIgzlGacG8XDJ689b2la7U3dcJEh2TNEXUblHlgCeWZ5OeNShiZxkZwPMIzcTXbaMjufVjXjOXk
uvGhJdaCrXkHXuv5KoUI7PGTy57ZwFX+07ReMFXR3dMitnrAkm+JYN3DBB7Qq1EOvw8pcc7WJi5M
wJzod/i73BCqWl+MdUk/CSIoD47y5gyZlMCBbzMgLJf1k3ZkTteynCY6FBa07qKNfRIPHizr21p0
OCFm2zMWfGL7MMchlsWJuUBxEwqMkd53eHzbhmDDQc7S8VxSrViZwqZmnO7aTVkEiio9CizuN837
KnewdcbItuvCUvX0eYP79Kq+LtiybmlUVPhNR4MU3aK1cyahOsc3bb6y8ci+I/oBKqPffyR8Ytxp
IpAhp067Pkks03X4IQ/9vKVztiXfc9hDivlp7jZxSoNU1YpGE4hmtUdcYuVMsAjzlEfcfeavWNu4
Y9hX/D4zYdHcnLZQ9TlO+BaYKtST5sWvVKcXsd9+712ICgtXDQwW9D6xjDVisBsW8Dd79ZewMB40
kzAOoQ8r4IVhrAVlnNKcuU9nwIG9wWW0dozIwOOZaX5fwSyC9lX/3vt4lPEIi53y1nSQNspzkVFp
3pxE7S1YZizsiO+1bhhoTqS7EvV/TDPcVcmlt53zxuUbX+Q/9jtiHpPvvYCnLLdjumds7erscC5C
m+z/xO3n14JkQQXl5LcyyPGqycqmt3H9Q+XM5aDVOXb5/27H3JeuCvnIRaMLZm+kV7L6ANEzVIBk
PbvosVb7+HE4j92HQV3HDGlthTGYvpX+yX1C4ZYNrfLhU7EodVWzlyYBGOrtakTqrEmK213jHSXL
ktvJKkWKf/QpWjVX9n78FU3gg5nLf8fdOERl2/LlbwrP9Ub1sR7qa93EbfLSatcGkFIDB6a4e6g/
IlXjyGfr35SLUwi8XAKEb112CvTn2/xGVMcdcBveQHLP6kEDxiEX5xIy4g1x8NXUnLYpEsCyD9yq
sAGCoHNAx3IXyKARzQHSE87e79JK5pWQd2EhGDWi1I01bHdN1dKaM6Z9vi+2LlXbfKHAU93SJeRx
MYKO3JJIJAPEvwydvU6bBaEVRRaHynwMFNugZNZCQerJxnUM1Ni/SiuJiA7JR02YVuBYZObv39uk
h/cNwpkuZJ59a+1zVb1UMAzgS0y6EoFbp2rvNmafdyyTz9KDlZd8tonGgi0JfnTf03/G5CEd4c/r
71SnuD7M/vUExF0I8nhs518Ty041113o61IDxpyOka4aqKlncaG7d/01MlQg3I7vBTH7J+UVeDcS
r50IcYvYYNCsP5y+s0vqfFh4WbZZsDGdz5TsCpTXshh0iiEvBxouK4UDvwvMF/LWaqqWGdRk2i44
B3ypt3V7UH6INLB0yfthssXvL6HPKw2xfBGYjsE0hQgk5Q9AMixrLfHFbcToqWpA22SkinVVuQR4
Vkc3mUyAUMXFLOeTcv6L5uB2TQFxChl7Hun86l2s1il8wbDDqXcQk9dDpzDK3ayTzX0htkQgYGLu
9KAjYfRmUJYUZSy4G6SKPPjaOnq2+ZT1Vg3RjD/4qUoQHgIsXUkHmfTqJXoZL/kakfnk6qlga3KR
N8TsH/eNyEGLY7e/sbK/PQ6L+lTgmXmgZEqSMC5/s6m7r2mutyITBpkbMnYSr5XK1oSeM81JBsym
NAoE4pRwnVmLdp8rdIfpfxCjk7KtwaNB8/BstW2kdOcxbhZrfbcxUp89qaCVn3NNApGKpJCdZq1/
LPxmn0eeAfl9Chwko6NZKOo2QnF9fTZre+2awWKlla4uOcWpMgmtCZtpSBXNp1fRL+44/La4GYrh
m8HW7jsxM08z+ty/34hWjJdN+1hO6GzcpYX5JaZSORuMnqxm9S9+sct71TEHcNaUwqacgERryt/a
uTpD+5UtBeQZxiptM1j6uGy7OdbxO3RQZV0uit1l0k4z+exJRgjkwm6IXh3eUxENCR2jQDppar0E
L254g+J+VbwbY4RI3Z6jm0fo1vsylUn2sxIDi7L2RJ9OtXBHRrYIhXyOv986xvGkezhdqLKq/vwm
P5n8z87z4N2VnEGSqchxIIXv7dsz+JrBcyxDBPLWZhpiV+Cq8Pextz+GgV6bU5BkZT76o1dx/eHs
6DPcFC0j+x7XKigHaUKT1m3nu/fA9043LO5umtJdQUPMebsVCPAACc/fualv3mKH6LMJACcogMeB
LV4v1zq6lrsJGAwUJF00DyEiBtZE9QF8Tb/TgIHJc5wom4NdbitolURbATnU8plpGey/5AjsywPz
kT1hua/c8daXzqXrPSXiR1mqiUOt3Ebq3wDfHh7ZK9hqMisGOgjWYb34BlfeqP0sceuWFCJiKLFH
AQmGwoCfgM0px8B1KgxtmGJFu7T8Yzs7Z32JriJQdiZ0bATVWLO5OKhBNreIEUsLkh5vvSInVTaG
fBgHoJ//PECIp71oP5XEU+ddjjONpkvYAHGL2w5QmyBqrUWxpyQlNbzhXWlLM2nyiRs5PywxXjgP
ZQkzRfuof1nvUPr/8O+ff8kFFEdmeKSLS/Hj6skdP8xuXLrI6ILcFY614QdnGKWS/qRIhiJlR99U
hln2XPRGLMsrqxYH2E3RYIpKo/ujgxfXXy4sTNy4jjvIsBN+r2fwSmWCLN0913QNm1M0ExN0fuER
sOPs3Y42Q42GjNoWDC7lZrJfvIlynBx6/eaVqsLkpV5mdSW/yeppebqQOiueUUXXf3pQg9RrOMqA
rBJFApSH1TjlYSoj1tVqb0eDCWdmzB0eljqzjom7RrRFY/DOi+6uML7mz2w00zUft/iEAcwNvkPE
3ezP3mb71Hx8CnuJXhCagiKq6dj1Qdka3iqrbDHzohpYIU7W31LlDgDfuNbD1ORcH012THrf53d9
G7mlTn68MmovE1zbaZ6qeh0euYUlf4CKnwb9cm/H6Jy5tyORIzOFIcjwgwQjPtVzGeu1bTONXsUU
pdLdvk8SSp5OnpiAhRHrt2xCUr/CYS44Dt0f+9hLH7wB/H4+1VHjzZBznWIxpJdot+uz/NPSoHdj
GzbSvUBkWOcxeNTnBvjhO8HrU3iNieiQuNUPBc8Sudi8YOOgEHxTUfdvx7hB/+ROIyZSe3PeWLde
E+/ePjfzZDpFzgG7Rp1rKBAOuMEjTIkbH/3Imy8QNw1SpEzqmrOf4hq9Oqq8fRDOVUyha6krmfYv
W3WnDdpGLi6QKmxn+OV0qZ4xfDG3aHPDsMlflETuhWRnw44PXPePSbRs9UfYKSXAagnXYTZ3vp35
saJLVaCbKdEnPhfVQZOiyXKcTGqEqYEe0cUwA2vyq7X6DSgrqEBPZB+fv3pNHzz6QAzQiiLvZBOU
LYBMe5VpA682FQ9zc4/T7WmvF0ZKMjK9EpZFvfn2uo9wUDdTO/4d0Ip88GAjanHUgCysmel7ebGf
fj1zImDgOc7K2SPEKPOBxkcNDhS9+cEPKJR1T63QMWp2wjsNcjrqE1/6o8YRS57+4nea/MvwdbQm
qTXTyXDA1vS+ee011FjjsSz7+YACJN47HG/gzLs67BeuxoT6LeVby20hpzz5Y1mgnt4ivkt5I2Wr
1Sq9G5Tfsuy36+3YEYX7fCvwmqe7t90k/PNX7uOCfk6Grd3nHEVsqI74+j/OKFom7/6JuLFNB1sW
2F/pkxJtwI+Pz59UQnmSCaEhfOWz/K2UMQrHPIEU3NsH5pwiXYlQpkPvhKlT6RoYeIIkTwtGIMKx
z8Gjk4w4eFrFCjinMpojEvel9Vup1nAPZpoIVonVrDdWemO+VIYpnYfoYLFGt1tMt3ZVEXZDbW5b
IqbfKmZnEt5mBwySOlMERbm0PN8tJ2cyc84HcaxywqKxFIqXNX2HVzKpMqLleNe1GO7NN4X4xxg6
mnXHO18fr+DwFNifNNXQuTMof1nScBfv9zU5msgmTOUjTLeAoaBC7wdlHdOz7SvL/ClwRSvnXqtR
TYD8rRegwXvR96+1740UQxwSzMDAePqfdrqykB2ZCJN2n7/CWVE8HUqQ1rZiA6W+cUcOFi730VVm
wQDFPavCi1AMt1A0G5anWglCKBnnxF8H1HHQf3ORRAjZrv5WPi9H9BzGkBfE6N7U9NgrwhsN8YUv
OEt4tGyQBUdQ3A4JE0lEJSShMrCtGHmFX5+OFeGycNypEwKkxiBH7G8AFqQf98tDq9e+8s0hL55K
RI3DQbegvz+loGyEsISUflMZBk16lmiEvsRMXVOkNV8JU7ekH4zCKDRAz8TLD2sgwkol6RZ/vR4l
QtVndeg9RNVjYpiZpt1Ih4HMSzGoi87FENeXW0LpM98XXOGcnMNqcyvZrxeD1CrUJH49UfKqnDxQ
+qpalmEcaLK9r1sTJ0kbjRc+DvcR9ed1XIKkfXJb54VDb9DVZMLWQT7TO30FvuUc99/2XOnMUS1q
x3OCg0uFSEaMm/2Lxng7kdEfGCrzjKrEvxcUCc7e4ttSPV5XLA/kptoHjWJCd7IKSlr/q1XBfhgw
1zd6WfrLlI9FKdROrkMUOXwJGy5TZsbTbotyooIAL9Q3/Ad7bwK30QyGJg8Rmgp+MNcTUoKuv7ZG
W7RJiz2tLk3jshQzFrN/hoeaDP0rqCH5Z8YRTwPLeOUTRB0JoNhM7E2sxQVyj8PmKBo+wp+Tmoxi
uWEOQfonWnUfhpFby2uclDzdzMjNHtTp3tfJxtE8zVo3ffOz7ivH0wmUh9JYECFWvZYbhMSenR1p
FFlTzBrTZkr/Vb/07X3+TZJzhzyFI1ac2CPM0VOpaY/ag7vv+6AuHptRueJ15y83EQTZkLl+TbMs
9e8nUTRBebY6ZR1asCJ/GRXl0OZakcm//iAWEVptROupWPPKwGy0yRPTRR8+W1g10moj1WP9Hh+W
9L109wyoP1EvJQ7mtiK8sc+qqmvRzthzbUHnZKAzvCj+nTRTk6HNXNbJk7uSQrILARk9ZVlePSV8
r6Q7m2vQJpEr0uyr69P+LV2chbRoH+BlTL4Co2XVwveJMHbIscSK571Sa28cXk/9Wb9eaGKsOcdF
LjKdT1oE74nKC9NE+pkX4++qrFWvz7PfjBkjbaGl7cVEso6r4FqOEol0AOZHncYXB33JZ4c91PdG
uM6/jwfKHLHA1mgDXr3QQLP0orpa4VVwuxhLED4ftYj8MYlYPJ62W6C4RrRRV0SldmymJYi5L++2
mtLwt8kSBaYGEVDc/G7yIy+KQqEVi4Pr83YCd7ObP1062S3xRWINlQdGgTTHxWPeBcbh8JaTt1tA
IyurhuNIx/TlSXFQHsZrhQHB6hOZsNqMzeeWIrmmAwi0Juc2gH9xrrpSVLsY5bD/iOSXbbZu1oai
RxvYTaYI12bh9bTxlDPd8oM4p9guQqzBaR9Wq7/Cl4JJZD9lJzqAt7Q8vTiYxO+iLOjUUsrKFE1+
8e0v/yU7d5vbj77YjO5RUdGhSXLLWk/3IVwZ5GwqFAwLo72HQj0GT1I0Ab/V0Wdr9g23Vygdhdpn
RDAaZvCQ/gUR4UnIPHMgz7yYRNdHaHYVRqXN1KZDjzBBJ30VXrqaYbaSs/O0NlUYWM7miJdOEFkt
rN9967u+SYVTsEU6OjwE2YnevwrQaeJ2RfnS8XlW158BVfonCUDK3qxA6ZDHW9icPjEZIIdyviFi
xq25CvNpZIhhBnPWyn3cwygfPYjXuUOuw1iH1ae0KttfpkS2Gx/+/HNsCppM5OOg+NTUT380deQM
pBxjI4QQUEwvAq7Dj+b/TeNjS9rAck+ooFZUNMnKYIlEqFefyZRfWZsvpwClhPVi4DyPqCFGiY0S
Zhta6dJjIhx2ljaHlesXYOIvSYQ+uHs9V7OkIttNtPqIZKlxjVzc7hkcF/G5einF2232ak6akOD/
1ywM2MNVb2R+pZcThn3hiH+XepDerjq6nvZsLh7WPSma83T+bTJ70mtYo4H9oQXNcnkE2qhKvf+A
tlb0ccFyJEFLjlRHuMDYJUWS1c036FvaZdWQOcQAgS+ps9ZHo/DuifF/yyDCN2YWp+WwBLn+vWYu
GzapcCVUUkhpNwvMWPKNxg0Z7LR9j702K0yk4Orrdggh3/UAIGF8jKez7z/2frbKmxGGRs3RsW+1
3vd+xjJCzeYX/Tz9FsD/b+mx1gEDgdoY4ale25adUtDgxxuRERgSO7w8bnbLMv6leD+MT3K/iIkl
kw6WlSBU5RGoodTmOa299lRzHp8e4N/WzR2tGQd6Kcp9iXu+MGODC7udIuZTx+3TeVgrVNai703M
2+ClXu8dEdb81LvdIlC7/3F9NOzg6aaR/WMq2VkZ9Qa+bnykxbOI4488CerHaoKeeHvr86zOiqYb
MLlF0/svtE93XAkdHDDdiHmg4jXStaROqeXVvg5d/gzYggQ2yZNh6qeNn2CFxgxyBweQCQ7+ugwv
aCidMpNKFqLkSN8sGddSylMKxlS+KxZqO8RFp8dohHaEXJ2WGgULFcEcTYxa8w5nSVfArCoxNjHy
7Q02XZ9DhDaIxJEH07SaPXZ13n0xJ1riWKUoEjsYxwYI7pmKdMyvkfLDnw82NcLhgL72MW5vMaXM
WeLNB9WOI8BJsAQPvvfL7AiXvj9adzOjEpPPqvFxVUUAq3mKwROPRqJU/NQPg4meJ06vxyNwDJHN
+BP1OJpWqQsn30NeeZtd4ta96booHPFhy3Qt7yQdpyo31SLxxa5X4ijMQbpNbQbWa3CbejzF6Znx
h3IkioI8B1BQFMSZG3MF9vprSYkMPm7367+N25jVwFxURKrKp4RYVbOMj0mctSY7S3Xbp5vmJyoc
gsdnkbob94wU2JrtgB3mFTi3vUjNT5rmbbzHZQuyJg0Xmg6qi/iKA7YvZtnrQmi3WCppZ9/tlpmd
ohO/9bhySMEu1Vvr/MsidkL/8Z5U2UWYVMN5A+VzFSF9YH9I/BcBTrkCLvoONluO+CjbGZRi6+ys
MEzDcCBEX0Q2W9GXokiQRM8UCWXGbihS7ZRSRo20f2DqzhSlmXB7muQ5nQCLgsK18k1YcbwG+It/
r/Q4SuB2cBs0P6YjtR6tRxmcbp9mqHx9SrtmxJklX14siL7uxXtxzjwATYwZAi9UvrXkh3dc0hXZ
R+woVx7wYoU9g8cWiHkSDb8rH4U0QHwveKYcTCYb97zqGvg4CiqUHYcYYE0jk6p7mObNi3peN8jh
gywEXGq0vT4NKQL+t+DmyKT4+OOpAhA1VFm8w+GZmPjHWu28jSGXSviy1n8xpUcebNcd59XlXBrD
GyGzkDqnF3KVf0CjtzsGi9Ek00VLhegfYmoDJbG5hiDbvf945bW29ihyFIT/ZfrNfcsq3QzX2cDK
brDDdKzzj39FLtG/5LST0mhAx1v3xFMZowu8Qy/jdBucnbG3ya0RowvUCmKsGQGC1TRSD3Scibl3
vHTqcx7GxV7TH2jwwDB6CVBN1DRylBVC6T+rbtzI6ghdYi/btvorMpBk4nVVkD9CiJm1J+HHezUU
JMNcZpjQdrddxhsgXK/8XTlA4CgRWTzrG+OTqTa/ZBfnZ+mjDH2PDQAFmWyCLdszyazym5ObLZXl
8vax90MFeLh/7HrLvV/7fSpveJwhjoXwn1rNVjHwPdiKdl5diRio/nu+IHWQJCxiom8b2WPpyXut
Vti5YQMcjJHc297byRiEtbHnE5kYf66VugolTDQhw1IL5alGnLM3NDbKK9LRNH9tvsZbGX+DG8Ly
riKg5d7zheHJvvUmV79V0XNopow7NdFimNeRFJULM4Lyt8HIfB26ty2RvX3sVo47AbMPpbG+DB5o
WfhaaOXVDO4c7vncaUAii7nCotQoI8Ephqplnbibwct2OHN/qLUSHrQ8v6hvGfBULYqCFDx8tSGS
pMDi+ToiOZvQ5TAdoCTvlmgbKcyZZOXohI78RWhlpkpjDrFa4Ha9xDgU8S/SX4HplqHuarss23GH
H5B+A8RpNHEUolV4C337MvPbxROLjs5xLHc8ntqCOmEp5kNrwOQGicmTDMUM+bDo9UKYpaM2e0bN
qQfhb/F3FH9iRce9apqCvn5vhfcvGWpO+a0KclGxzC+RejM0dqD/DtrBTDBk6ytFxM3Vv7kYsI97
YSwWo6VNzH+Pa4vKUB1aT2ZDYLpYYs9vxrH49NXbEXTilXbp3F/MJhaZjlMXgE/IY33CXPYNaMed
qnIZs1yTdp/nd1isdYAnuPEucBdCh9U1lmv1DwG9ueTT47A0b6TQ20gfDp+OS1GRyLyQrxyCe0na
hOwtG1I2Ujq5sUMQSMaqXk/S9qB6spCEp0VzJ38nHiwWernVn5Jd9jPxlaNDPdL1orxp1rnbfMI6
5nDbhE2ppirAg2xs2/AaTdpJP/RXf9oPShU0vO8MvJxMktCU4PTSQe0teZwJwbkMvcwTlmlaGp7I
gMBNWQwed/4cBRfj9Ov5nm1nyMav0gSlY81o20OykmwR/ZFM3nUwcnu5S1INVetjx9vV4RWksv+Q
CptCUCSOFOWwlZn8NE3Zs3OizdoX5E2MWocU3Dz1VBbVPZmjP/nxmb/T5AG99IuIVZHaXmukeF4H
YWRKguyLlIcZ4O4ZaeEW7qmvSpXrl2bTuREY/7XBqqEtJUJU8c07zNKfRDgGPY6VcsGEojful6UX
juXD+k4sKCDMYGD9G/xANzXyExhgjhSjKcxzx2momBLkljJ6N0na5WKuIbtEchsXtCd90RhBpbQ3
/6FntqxkooITHWN5B7teqse4qXRBDg1T4dJCHvEUI+OKcfPobzM+mihh7VMilOCgjqhdT2mOIabp
dO9bQ6rIzroBCyVDK4lhp05mHwfPqMiP4/Xu6Bqw19w4Wc+3GOOCzvWjuf6EHyq52J8waCJiyJkV
lrROzk8KTwgfdSdkrKezZF8tYEYaEFXQl/DqUieVq9lxAwkZ7j/luMJZaeTAbP0cT/fMe6SehpAe
LtGh95FRJc3gvtpNKcaOjG+qt/BrLN/JjG7xPQ/A3JzjYrW4TTxqiuQAOeyJ1f8R7hymejfcUb3y
L91yiESKFwc16esj6hXcDEwaGVm4+zhQHh0j2QikEEe3zQt3X40kCXRBrrDpW4q9myaq62JjAZ4d
tsd4t7bAfqc4buPlJohyWFF96q9hREWf3YVbJ9dlMf0l/L+/ZUkYDT/oIKawrOfqzaTOoD47UxSY
cX/xQQs6QWu3CJeE9Q+mvN61iY5xV50SOoJnQD/zbZO96dFOUF7D9p0cDBTU/y6AiCNlAX9TlWIA
jQINbK2ccwNPDPq6GubcckkJMwRtUpaax2ZHLHSocBkjdk7nlVndyMBEZf7x6MFjrFALJTJJsuiB
Xzhu9N6dQ6o9P1EF9JScQks+Eo/6wRYEkJYMmj2T97Z6dmZGSW0vkY6zUpoaMfcVICk9mLA7hvdn
9Af11TXJcqsjLxklHlgVAWzV+qY7AADh5uUTmAyZGSQutCoSCfTkfYgpiyTlf3mxyGlu+xZ7/He4
1LNZCnGLZT+LS4jwEqWlluk2JV03hJJ5iRJKXvUdWBggr5H/Wgv1kL1BHUEKVSsEHsQZXkudws6L
nY9iUCVMP/lcjLEE6M/cFudN4heAXL6med8Yb2W6XIkudzj2OuIdydK7mNU2Ce52fkadmQ5Mvm+K
HuZu03QyNCWK1EhPpnWZOetc/FeU3b0vsaBYJ8QvexDmeMvcDfMc+2WwrkKp/+GyOnKF9qDfwH89
Zu1TnmfJg6RNcoSY/abQ3SaaxNVoXF0eOu6yfZUkCV7nKU34sYfKXKuLIPGdFfvQ7UeiFx+S6N5v
79cN2ONHNDt+9bD0hvQnB/Qb10pwcVGRRTN7mm9X4xZJaVahToCzy9kMXXI4x8DcuPZ+K4LJsGeR
MvEth0oSr11T5xcbqiYB1gd0/eHizqEdbcX4jQOQSK5Kfn0Xu4WJfY0FUAE2s1MrowLVs16GpgiS
Mh3tczq2D7DdFJLO09mOqY910cCpJA1aihkESJYmR2xl8Hjpq3dGX9moBPuUj0HSozAOO1c55N/t
rUBr6JDV5uQCWY37OmbFEtqFqvDLf7oHng0np11svwLyGPgWfk1PhIalih/DkKGATODUskSeQ3Zj
R6mChG/dq6iGDgXGQJ6NPnl/DNnehBTtaWEL1Wze+PUTuHxjFvX0LxXCBgBvLDD+gn7OTm1me6bN
x8+SKLG2MXYhAT3Uy625FHpyFffXWOrL+/wKHnE7iG50aorSRgOvbCD0pcZSgCCeY42erMcieNDA
35UrllI41ASgULzGpB5g1J9WKwJ7s+79V0xvIjLR7BUwPVXcwZhyN1Y5ZtP8ATAj/Xs3qW+EA/PK
bbk+rvwlhrW9NzyL5/BC030GxmJmDiaZ3Cjcxs+bybc3OMxQGpBY9n1UUTfHOxXlyH+S+oG/4o11
2eEVEhEq03EqkQcerbvNLUwfRSf29vOwZ5WR+UQlR+QWtDljRg0Vv8leWESFg09CisAMcL6d73uL
e5rtSGix6JJh28d47S213e8no4sFYgtaRYYy3Tnf/5DN7/KdS+65o2jHGjch4jozXwrTHfjXmJh5
GWPbl8fUvr17yo/0LsLhQkWDguB6o/e95aqIpszGHXzjyyav+cLiwJADsEC/CsN97JEBgjoAChcW
mX9k0stwvmXsthJzot5Sec8qAXVE43cyrgEcdhn2MMyWgWAT1+YQmK54DwNMhAmkMMrBoCyYGUqf
9DYl0hDg+Qvm6Yy8WRnBmSXK6dWegcoY1MZZbB6xCJmAeM03OKLeDEzpbvDks4oCZCIF2wgHj24Z
V/2UrE36sqBFYPe0z6dvrbetDrt1fubLSEyqBSaLD31RBdinGIkaiSRDjaIulfW/pFHghX/FOkkg
JU7YmcXvP8wuLWy+GhozLG0CJw+XwPMdcqaHx6bP8N6wn9VQP7vv1Ua7XLi0HBd57A+MuoX1uqos
OLlt9lNCjdZ6QjOiII58JQSpVuMfrE/BAUsmCYid6MIvOeZyOA26DXEPiFXvosqUbsKMEuYRyzgY
XQN25j/pmVL9zOpdkCj+diTPaHo5K5qQn8l5j/19lvps+pqudi0s2+UXqzR+OJmM5fmBAIisOjnN
4ABbR5Da/iga8sNjfWZ219+imSoWQdt31iWanrJ7d8hwVSmVhA8n5wO2QvI3hGZq/n9RGG8CcIxJ
2fpskvD3BcumijUWLszd0JcjZaHG4qz++CRG1B7+UQOgLJiq2hAVkxxuijJUDKoYXRImMVP5kOXe
uGTkJlfrs0yIMZtOfBsox3Zc4hXggzucxyhOSMZsJSAud5ktEjaB/cNK6DJuOozDsNcrjyeshUEZ
GcK97hIvp76hNoC1NMwmdcBJQDcCOv6ZQtsvZlNimU5AdnkIMuv34d08lyxkGyryThggAkob/lwi
dbz23P6yDRBeKzRJp4BqkYo5HIX8TRyWgzgydpOlS/d4CgnJ9Z+5BL2CD+n5Y962s/M5cJamWJyN
TrVBpe8JxbvDcFVoa8byu8apTLAo+kw3WuXfrIfAio2PuRwfKm9vIwlV+L2+5XuQVvCE20NVmMxm
YQaAvFRD0HaNnDUTcGJpktSzOYNBG539+hmbjQn8Mlz5i8Bf16xDK5U5lQW1yJqziYLAXwOXLp6N
kgEmbJHn+21FpO3w3NueFFAIHGjtfsaZXZAugLVCszDiCb0/L6PT2o5i0NZUFHciRF/0H4mHyF8n
kEyNgZFT0dSdW9byziqLcLPC09P3JRqlunDACyB4z2om7rshYsUenUDsEPRPfZwUsI+TDirQwq0F
j127m8tn/D+dlyRi4n8zOmmeIqM1uCCchiAPPr9nLCo/+R3+HI8yONF73d5JTujEwLwmAT/VlDa2
pKvFBk6R5sblmF9z4mdLQIKeoppl25wVStx40OaC+S9vOhvUWMrYG317pqH84ijCH3zg60NAJMS+
Rkl1ZYnEfVKI4nt8oAGEE3V/p56KowejZXuHB2sS+vCsodvUHlIe2Vk5CrgQpCQFpt15zG+E4iD6
DwtrpeDniBuPezgNhI68cvhrBvhNdM2/UWpQmvbKZazawjHqgW9+JLwXi+5RvET28kcpXLidw3cN
4B4cXbaQuZmc/LOh71kewumHAzxOwx2HxDWQWpWN9srnDSLCvnE0x/fRYuVLLHF2hsv7bkVdfyhr
chJrhrXaz9Iyt8JHv4ZD7KyQ0r98EMlIXiKbzMqnv3+qpOQIQ5WcmKIS7IH/3yXeL0S9bngJbFwS
SXNMEjyJJGLyYgeDCaP1nMwSNGJ6Ycwy/ZpXVzaJreW9qqXYGekQNBGoc056JQI5lTOV2p/Y9A94
vkhCO3E0bmp9art0j0gEE1wpJvRRT4Q9gJ9crxEIWNM3Mw89KBuBl1J4LAEyioLxZUkNpsiEI1a3
zgXTEtzLetrwJI+00q59dPz+u9vlp5fOZGp9IPv1eoyINEGu9Mn/I6PzgppF/IlkTgX7MMwpreRp
oMo0BrrLesAyUQXaBaK6p7rncml4NaLFgZnxRP3wdjEdEklMlrqjrhNWBva0qw6Kg+0r0+Dnjhp8
Sl7YcjaywZ5x2Qng8EI0mm+zWF0pQwrt8nESTprF3xKQpCKM53rI8k4GLLmKXZJjgDS2MVepvdyK
qFnPI+31D/PZ5Kyt8MlkFLd729vfm6J3+39ic7uN4ZcQkY0xdcwCmt4aF132m+G0idty97xgjl30
XBqgjgOf6meCrIRcamDTlZQlA4hIZf8yCnj9AFiz3SlpR+NMCx6lET/Ct2Czb1v5d5rR0m1xL7MA
n2CF2Sr3U4fBjyTSRdU8o8KTK2YqyoD1k3gAQz0oKkSWChAd1DPWv5aXfzW+yfFqFSAVJtzBGSPn
sQXE1GUzecLhkCgqFvD14ngHrbzK5TtpTVRCxoI+mw5PqldIOyaJQTltzybLYuQqBKgCvpGrBeQT
3qeuEZfSGE1LiKegEAJyqyySFyk8FsqHXf4S7lsX++huM0fKhKIKziBZ9vGuve+cBsP/Euq2YHNa
Gt2WvVNLDfgbfLZ7zoW6+wbSaFfZ0r45z8nBYTlW3B7//kDxSY05Q/mwvE3+afd9IpHqg3grHNH5
Sqp6i5rCjubsdp/yM6TGBOKyl3m8T87e8byVvdoTjSqdPsBesB+H/FDTDdzwslU/qPp/UaTZKo0G
rLdQqB/lt1hhKTGXtQ1nledly8LjtAUSyuSagcJjHQCvNLhiq0tJ0a8yeo+/siSVn87muEHoS/c4
FYJVFG9Hwfu77b/lRjSufI+HPlOVXtAswLwXyfK0Ai+4VagmSk2NMZQDsm5s9Lon8CYJWt+mhQ6I
1Ck+0EFB6Sw9v2MbPzgFPYzQ1162yvKm6ZZ2ZB2COehzI2jjFgr7YBxYNpamyvk7x9/7fmoj84mw
BvJcm9++4pT0HQ36eSW7F156ZYUWCJF6v/xrLBaCbCtWhxKW2qRYZlf0c1vJwA7jDfCLMacPzTV9
CJOR/X8q0NCgl1cyvTxeQpzCvC8j/O1urDffUv8cNVa0t7yy6Zojp9UcUy/L2vcQcGQFWO1hEbqH
13gB9RJVQDJXmzDQB5dB5W8th0p0HmJBGTu+mCH7iOBtETi2NKqwF/yo+TXvNmpvOyPraHksmx9q
q3Ouazxg3oA9et9wEKIE/eXQWBVv6tkjSHmQWTE/0HaePkpRBD7uS4xBfPn/jYZoTEzFdxQujsqW
s9WOrWIO1n1+6uuC+gdljxmVK0tKNaXZKkyF+kvnmII2VrXkc1O8I4hvkMaadoD0Lo/Y3owjFut5
LG+5o3WVR4CK0ZOclZraDQ3ZdFJecMFdDcgrIgexMGU/KBMx70AC6v/cIRacbMud29V+SLQJOjD1
GniiJzsiEVvEOw2rBLz/nYgNWO1HWGpaWjoA+l7CvBjBjndHb18Au6Ks27FByR2kNpeVpehBhOEj
JvmSQ6brX9leF+KMdEoK0g/sHEdnLly85B6qfIEOGx3IhSpBWREiYY97f676Uxa+l97zf30AFsQq
OPVByPfiTZ+tRDOFMY8RaTDfnDSBbEGjvskOGcwsqdtC4oq+3stkj5axFzmPfmDRgu/q1kVPFAfF
O2EFOG5EFPK4z+aGWmzt1uYGccGVSM+mq/sI2riY+arFDauOCHWVuIGauz+54KSVGgEvK4U23SLo
VZrIe40IULBG2Lg8NmTw7B7a05y5tasWpxQ0c6x6N0T6x/NjkIPpSxMw805czjpxWHvRAgVDiRjs
u2r0SvSLUOqCdHdkhXJXQZRrahclCAaohpGtphnMdDkkq/oaBUO5yC625QbY6cFH4qok0x4UqciV
9eyJJvVcxHbRovDBaEbDIIiUXR7sNTGUFJAwCv5be8705RjW+zl6A5k+A50IQi95JtWBH1PjqbTs
oV/9QS71KH/5nkuhsPJ3V9dRKfUbCummqM0yPIM6WjwHm6yoEwFp9kh5EIwDDhH9hYHH8JfcQDtU
JKjmwY7XvzFZra3FPWQlD/XiTKNTeijCCpV1X/rFFsLkytA8uM+JP+B+0Gw6fAupIT3vIm6cxoer
2Drzr0cfHEeaDrdvoZURRW9HEPPLMXhOQSbbkN/XI+cZ9HP+YL96tJXtRWKGIa5XgMFEW7kkHLKl
5N2DRyfs5Cq4bTpDg0ZheXsDhhVer0KA0GmfrWxDtIz4hb7g8Jc6tBhx/3fMZ5RdHVowZSwt8Ts9
JU5em2LWJgzZ8IZ7wY6T7hKKDb3oqKqsA568DgHDzDubCVNdtgA3akQOKR74PRDZ+PATD29DsJdw
9o0SNzdbhH75MnMX0hnOv91JbRseURuyDx+YYr991b7WvVzXVxIozEZd51uHyy9aaHKwqgBy/JMt
K66tdpbkK9w2WXcf3K0xl2wLzMlJd33tgFtSiBYdK4cPattWbBsnd6aWE3TXNfApgm0KFOj/yUeD
h22sSGFWWySUWOLUh3ispFHGvpKW1RXvreAm0ouuiv8650uYj2VWp0vSAMGfUY5HReij/+oGZOgT
W3h67MOXM22X+gbdqE3NVzXv5XwoMxuBDfHzO3lZsMGWh4aUrKrVZwzsj71CNJMYPrzOlBkdoq7m
GWbbsqTexfodZ86l4pAnypjIdAyneKE49NxWXLDaXVGTrNJZvAV5VOjE6aFUA08V+Oi4lLBz38Ez
Gcw3XiU7GoVAPJ3QAOBZy8mW0MMxsEpR8et2TLwmOhkif2+mTi9f2o1c2UFHTx2Fr+2VROhvv39Y
WHZS9nvmj2nkyP7npCOyCjvtcSo8pi3rM5KYG9WtAqAG+E9sYqkQ3E6crVcWZ7kmbHmBL+KdQd0p
oJJ8cJQmyDtxmeK5od5rGL7dAVyexWOuwmH7bcfvCTQgqs7gpgIYmI/lc3wyBQ2vXL79rRlhP7cg
k4/3wQgcENTMjLPmRr9kVDvmS8zs9ea/j60r23E2oRPnpgg58kSTrIP7oCM3BbjuYAAd4PANQxJf
vGmpbu83msjFF7ipSH/OKfPT7AFnaE5JKsF9mN6PsqlA+CN18Wn9Z53244Y3EjetEYQ6TyarJJYe
GLt6julWKKvStBkwP0mxLyiLh/ITjkIX7JaKvHJozBoOMADRZTUy3WCjr12pbri2eQfyxR6o8LJ/
nZ2jcrh5rYe+q1UBPX5X1YUoPEUnVUNUx/vJvbPdKrE7eH4+cXWVrTv79RFTuI6s0R2LDllcAWhn
YZsa6q3NzDrPtNm/lljw+rLV15bLvvbcQHM9MCGkx/5IbhB5UST31mWKEl1o/6dT8leZDMWHuOSw
Zz7SLgSzYRKWJDZmYI3q5TdgKJqLFGa/eDpOvQvcl+rbLiGVqczw5o7U/liWWT7t/y+0J83+2rCL
wjX+5iYMCybiXQKFICWwlvCvLF7cCGSyn1YH99X78PmdF6Rn2Jh8XolbG6R6/2m6+/QdF1cdApn8
gluTlE9qo1/TAYrl77HwQreX/6kYmpLhU7/vKyhUoeKWngaQ6TNtLX4YWVD/eO8MmH1OGDwuqj0v
rVVmsG0qyjmSVIvwhLci8jkfc+J3BTlDP+2LsGprzJcUgYKORK/BBRinuHVkrQPntWHoxsWqT3Jj
uMBE9i8gs1tOf4qDaXGli0x5DZjp7ynttdIwOaVdJ7BjccuWqUdnYBBnny6J46ZPTWKInKpSzQI9
etRN86U+ybwGwNgMaU9sMZUPIoRhipwyzKyIoXEpHxmub2KzyZIPT/pRFTu5XBxNKMqXHhO9WJQo
j9eb72bIdX0AP5C57xRAWKhPQMK+0doIHBmQ++EIgJSZh/6/Ef5c9HTu6xNSlz0b1k3O9juBdb7s
xFZtPY9eHWN5ve+Mh0jEThq0xGGjIZfadxjZv0lE5ahIOfPk138qMSNC0H8zYOEX0PIhc2Oh2bsc
yHq+E9jXNrP2FJznoJMhArrkKGSsuaHuowANEAxRJmg9B/wKTs1w7WmbYzBAcHLQeh3P5PO4nXll
KgA5UlK1lzEqpkmG46P6DRLkdSYsW3ZkcnUwHEEl92Fq8lMk7MUmPdc/STRqNnqpD8DVon+gHmCO
fqp6mMmPmGPYiFfrKq47iQwmyCEvwaD6X2dFxoABAqErOUDMBKFssEpLY4TU7681e4uj5Kxeiai9
iYGbfGm4nkBEPyC3BqLJ6ZD1e6Fl9M/3unX/H0y4tdthqG6H338v7W7pHA4PSguyz2q1J1t3/Ff1
1oOUdpgH8OCV+/FmeAfYVNF+YHsI8YeFxz4KsDvKjZfC4AjAQ/58/3k/4NVj9/UwbJTrQusp2IML
75lnwh6tm+aUCOEQg2QVGZ/ZfM0ySeBES09gcAdz7N9NhMsCHRtuKsc+lyysoygOfweJIwgJe9UQ
AHNUGHxPfB3gotFjNwFudtNocRO2KedYIESg8Ztb9i7eUOTxn8J4KyVDGe2kwghUHKB+pW0KmTs9
dRIaeDqLhWzhFfjFWiOOIm+Nm/rj5T7D+jzX97nAC//U
`protect end_protected
